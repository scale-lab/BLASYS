module c5315(G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,
  G59,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,
  G78,G79,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,
  G97,G98,G99,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,
  G113,G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G124,G125,G126,G127,
  G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,G141,G142,
  G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,
  G158,G159,G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,
  G173,G174,G175,G176,G177,G178,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,G5201,G5202,G5203,G5204,
  G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,
  G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,
  G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
  G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,
  G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,
  G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,
  G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,
  G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
  G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,
  G5313,G5314,G5315);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,
  G59,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,
  G78,G79,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,
  G97,G98,G99,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,
  G113,G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G124,G125,G126,G127,
  G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,G141,G142,
  G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,
  G158,G159,G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,
  G173,G174,G175,G176,G177,G178;
output G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,G5201,G5202,G5203,G5204,
  G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,
  G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,
  G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
  G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,
  G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,
  G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,
  G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,
  G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
  G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,
  G5313,G5314,G5315;

  wire G632,G633,G634,G647,G659,G671,G684,G685,G686,G687,G688,G689,G690,G694,
    G706,G718,G730,G742,G746,G749,G752,G756,G768,G780,G792,G804,G813,G825,G836,
    G848,G860,G872,G884,G896,G908,G911,G914,G917,G920,G923,G926,G929,G932,G935,
    G938,G941,G944,G947,G950,G953,G956,G963,G970,G976,G980,G983,G993,G996,G999,
    G1002,G1005,G1008,G1011,G1014,G1017,G1020,G1023,G1026,G1029,G1032,G1035,
    G1038,G1041,G1044,G1047,G1050,G1053,G1060,G1067,G1070,G1075,G1081,G1084,
    G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,G1117,G1120,
    G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,G1162,G1172,
    G1184,G1196,G1208,G1214,G1218,G1230,G1242,G1245,G1248,G1256,G1264,G1272,
    G1280,G1287,G1294,G1301,G1308,G1311,G1314,G1317,G1320,G1323,G1326,G1329,
    G1332,G1335,G1338,G1341,G1344,G1347,G1350,G1353,G1356,G1359,G1362,G1365,
    G1368,G1371,G1374,G1377,G1380,G1383,G1386,G1389,G1392,G1395,G1398,G1401,
    G1404,G1407,G1410,G1413,G1416,G1419,G1422,G1425,G1428,G1431,G1434,G1437,
    G1440,G1443,G1446,G1449,G1452,G1455,G1458,G1459,G1460,G1461,G1462,G1463,
    G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,
    G1476,G1477,G1478,G1479,G1480,G1481,G1482,G1483,G1484,G1485,G1486,G1487,
    G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,
    G1500,G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,
    G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,G1526,G1537,G1548,
    G1554,G1565,G1576,G1577,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,
    G1590,G1591,G1592,G1593,G1594,G1595,G1601,G1612,G1623,G1629,G1640,G1651,
    G1652,G1663,G1674,G1685,G1696,G1697,G1698,G1699,G1700,G1701,G1702,G1703,
    G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,
    G1716,G1717,G1718,G1719,G1720,G1721,G1722,G1723,G1724,G1725,G1726,G1727,
    G1728,G1734,G1740,G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,
    G1750,G1755,G1764,G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,G1782,
    G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,
    G1795,G1796,G1797,G1798,G1799,G1800,G1801,G1802,G1803,G1804,G1805,G1806,
    G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1821,G1827,G1828,
    G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1842,G1843,G1844,
    G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,
    G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,
    G1869,G1870,G1871,G1872,G1873,G1876,G1879,G1880,G1883,G1886,G1887,G1888,
    G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
    G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1911,G1914,G1925,G1936,
    G1941,G1944,G1945,G1946,G1947,G1948,G1959,G1970,G1981,G1992,G2003,G2014,
    G2015,G2016,G2017,G2018,G2019,G2020,G2031,G2042,G2053,G2064,G2067,G2068,
    G2069,G2070,G2071,G2072,G2073,G2076,G2077,G2078,G2079,G2080,G2081,G2082,
    G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,
    G2095,G2096,G2097,G2098,G2099,G2100,G2101,G2102,G2103,G2104,G2105,G2108,
    G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
    G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,
    G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143,G2144,
    G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,
    G2157,G2158,G2159,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,
    G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
    G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,
    G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,G2201,G2202,G2203,G2204,
    G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,
    G2217,G2218,G2219,G2220,G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,
    G2229,G2230,G2231,G2240,G2241,G2242,G2243,G2244,G2245,G2248,G2249,G2250,
    G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,G2261,G2262,
    G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2277,G2278,G2279,
    G2280,G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,
    G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,G2301,G2302,G2303,
    G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2314,G2318,G2319,G2320,G2321,
    G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2332,G2336,G2339,G2340,G2341,
    G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2352,G2355,G2358,G2361,
    G2362,G2363,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,
    G2376,G2377,G2378,G2379,G2386,G2392,G2398,G2404,G2410,G2418,G2424,G2430,
    G2436,G2437,G2438,G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2454,
    G2460,G2466,G2472,G2480,G2486,G2492,G2499,G2500,G2501,G2502,G2503,G2504,
    G2505,G2506,G2507,G2508,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2520,
    G2523,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,
    G2537,G2538,G2539,G2540,G2543,G2547,G2550,G2553,G2556,G2559,G2562,G2565,
    G2568,G2571,G2574,G2577,G2580,G2583,G2586,G2589,G2590,G2591,G2592,G2593,
    G2596,G2599,G2600,G2601,G2602,G2603,G2606,G2609,G2612,G2615,G2618,G2621,
    G2624,G2625,G2626,G2629,G2632,G2635,G2638,G2641,G2644,G2647,G2650,G2653,
    G2656,G2659,G2662,G2663,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,
    G2674,G2675,G2679,G2685,G2692,G2693,G2696,G2700,G2705,G2711,G2715,G2720,
    G2726,G2727,G2731,G2737,G2744,G2752,G2759,G2770,G2774,G2780,G2787,G2788,
    G2792,G2797,G2804,G2810,G2817,G2828,G2832,G2837,G2843,G2844,G2850,G2857,
    G2865,G2872,G2875,G2876,G2877,G2878,G2879,G2883,G2887,G2888,G2891,G2894,
    G2897,G2900,G2903,G2906,G2909,G2912,G2915,G2918,G2921,G2924,G2927,G2930,
    G2933,G2936,G2939,G2942,G2945,G2948,G2951,G2954,G2957,G2960,G2963,G2966,
    G2969,G2972,G2975,G2978,G2981,G2984,G2987,G2990,G2993,G2996,G2999,G3002,
    G3005,G3008,G3011,G3014,G3017,G3020,G3023,G3026,G3029,G3032,G3035,G3038,
    G3039,G3040,G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,
    G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,G3063,G3064,
    G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,
    G3077,G3078,G3079,G3080,G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,
    G3089,G3090,G3091,G3092,G3093,G3094,G3097,G3098,G3099,G3100,G3101,G3102,
    G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,
    G3115,G3116,G3117,G3118,G3119,G3120,G3121,G3122,G3123,G3124,G3125,G3126,
    G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,
    G3139,G3140,G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,
    G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,G3161,G3162,
    G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,
    G3175,G3176,G3177,G3178,G3179,G3180,G3181,G3182,G3183,G3184,G3185,G3186,
    G3187,G3188,G3189,G3190,G3191,G3192,G3195,G3196,G3197,G3198,G3199,G3202,
    G3203,G3204,G3205,G3206,G3207,G3208,G3211,G3214,G3215,G3218,G3219,G3222,
    G3225,G3228,G3231,G3234,G3237,G3240,G3241,G3244,G3247,G3250,G3253,G3256,
    G3259,G3262,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,
    G3275,G3276,G3277,G3280,G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,
    G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
    G3301,G3302,G3303,G3313,G3314,G3315,G3316,G3317,G3331,G3332,G3333,G3334,
    G3335,G3336,G3337,G3338,G3339,G3340,G3341,G3342,G3343,G3344,G3348,G3351,
    G3355,G3358,G3359,G3360,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,
    G3371,G3374,G3377,G3380,G3383,G3386,G3393,G3404,G3415,G3421,G3428,G3438,
    G3449,G3459,G3466,G3467,G3474,G3485,G3495,G3503,G3517,G3533,G3546,G3552,
    G3559,G3570,G3576,G3583,G3594,G3604,G3605,G3606,G3607,G3608,G3609,G3610,
    G3611,G3621,G3629,G3645,G3658,G3664,G3665,G3666,G3670,G3674,G3677,G3681,
    G3685,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3700,
    G3703,G3706,G3709,G3710,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
    G3723,G3726,G3729,G3732,G3735,G3738,G3739,G3742,G3745,G3748,G3751,G3752,
    G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,G3761,G3762,G3763,G3764,
    G3765,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3779,G3780,
    G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,
    G3793,G3796,G3797,G3798,G3799,G3800,G3801,G3802,G3805,G3806,G3807,G3808,
    G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
    G3821,G3822,G3823,G3824,G3825,G3828,G3829,G3830,G3831,G3832,G3833,G3834,
    G3837,G3838,G3839,G3840,G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,
    G3849,G3852,G3855,G3856,G3857,G3858,G3859,G3862,G3863,G3864,G3865,G3866,
    G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,
    G3879,G3882,G3885,G3888,G3891,G3894,G3897,G3900,G3903,G3904,G3905,G3906,
    G3909,G3912,G3915,G3918,G3921,G3924,G3927,G3930,G3933,G3936,G3939,G3942,
    G3945,G3948,G3951,G3954,G3957,G3960,G3963,G3966,G3969,G3972,G3975,G3978,
    G3981,G3984,G3987,G3990,G3993,G3996,G3999,G4002,G4005,G4008,G4011,G4014,
    G4017,G4020,G4023,G4026,G4029,G4032,G4035,G4038,G4039,G4040,G4041,G4042,
    G4043,G4044,G4045,G4046,G4047,G4048,G4051,G4054,G4058,G4061,G4064,G4065,
    G4068,G4072,G4075,G4076,G4077,G4080,G4081,G4082,G4083,G4084,G4085,G4086,
    G4087,G4088,G4089,G4092,G4095,G4098,G4101,G4104,G4107,G4110,G4113,G4116,
    G4119,G4122,G4125,G4128,G4131,G4134,G4137,G4140,G4143,G4146,G4149,G4152,
    G4155,G4158,G4161,G4164,G4167,G4170,G4173,G4174,G4175,G4176,G4177,G4180,
    G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,
    G4195,G4196,G4197,G4198,G4199,G4200,G4201,G4202,G4203,G4204,G4205,G4206,
    G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,
    G4219,G4220,G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4230,G4231,G4232,
    G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,G4241,G4242,G4243,G4244,
    G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4257,G4260,
    G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,
    G4273,G4274,G4275,G4276,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,
    G4290,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,G4301,G4302,G4303,
    G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4319,G4320,G4321,G4322,
    G4323,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4339,G4340,G4343,
    G4344,G4345,G4346,G4349,G4350,G4351,G4352,G4355,G4356,G4359,G4360,G4363,
    G4364,G4367,G4368,G4369,G4370,G4371,G4374,G4375,G4376,G4377,G4378,G4381,
    G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,
    G4394,G4395,G4396,G4397,G4398,G4399,G4400,G4403,G4404,G4405,G4406,G4407,
    G4408,G4409,G4413,G4414,G4415,G4416,G4417,G4420,G4423,G4424,G4425,G4426,
    G4427,G4428,G4429,G4430,G4431,G4432,G4437,G4440,G4443,G4446,G4449,G4450,
    G4453,G4454,G4455,G4456,G4457,G4458,G4463,G4466,G4469,G4472,G4473,G4476,
    G4477,G4478,G4479,G4480,G4483,G4484,G4487,G4488,G4489,G4490,G4491,G4492,
    G4493,G4494,G4497,G4498,G4501,G4504,G4507,G4508,G4509,G4510,G4511,G4512,
    G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,G4521,G4522,G4523,G4524,
    G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,
    G4537,G4538,G4539,G4540,G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,
    G4549,G4550,G4551,G4552,G4553,G4554,G4560,G4561,G4562,G4568,G4569,G4570,
    G4571,G4572,G4573,G4576,G4579,G4580,G4581,G4582,G4583,G4586,G4589,G4592,
    G4593,G4594,G4597,G4600,G4603,G4606,G4613,G4616,G4619,G4622,G4623,G4624,
    G4630,G4636,G4642,G4648,G4654,G4655,G4658,G4664,G4670,G4671,G4672,G4673,
    G4674,G4675,G4676,G4677,G4678,G4679,G4680,G4681,G4684,G4687,G4690,G4691,
    G4692,G4693,G4694,G4697,G4700,G4701,G4702,G4703,G4704,G4705,G4706,G4709,
    G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,G4721,
    G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,
    G4734,G4735,G4736,G4737,G4738,G4739,G4740,G4741,G4742,G4743,G4744,G4745,
    G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,
    G4758,G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,
    G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,G4786,G4792,G4798,
    G4804,G4810,G4816,G4822,G4828,G4831,G4834,G4835,G4836,G4837,G4838,G4841,
    G4844,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,
    G4858,G4859,G4860,G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,
    G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,G4881,
    G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4895,
    G4898,G4899,G4900,G4901,G4902,G4903,G4904,G4907,G4908,G4909,G4910,G4911,
    G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,G4923,G4926,G4927,
    G4928,G4929,G4930,G4933,G4936,G4939,G4940,G4941,G4942,G4943,G4944,G4945,
    G4946,G4947,G4948,G4951,G4954,G4955,G4956,G4957,G4958,G4959,G4960,G4963,
    G4964,G4965,G4966,G4967,G4968,G4971,G4974,G4975,G4976,G4977,G4978,G4981,
    G4984,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4999,
    G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5011,G5012,G5013,G5014,G5015,
    G5016,G5019,G5022,G5023,G5024,G5025,G5026,G5029,G5032,G5035,G5036,G5037,
    G5038,G5039,G5040,G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5051,
    G5054,G5055,G5056,G5059,G5060,G5061,G5062,G5063,G5064,G5067,G5070,G5073,
    G5076,G5077,G5078,G5079,G5080,G5083,G5084,G5085,G5086,G5087,G5088,G5089,
    G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5101,G5104,G5107,
    G5108,G5111,G5114,G5115,G5116,G5117,G5118,G5119,G5120,G5121,G5122,G5123,
    G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,
    G5138,G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5150,G5153,G5154,G5155,
    G5156,G5157,G5158,G5159,G5162,G5165,G5166,G5167,G5168,G5169,G5172,G5175,
    G5178,G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,
    G5192;

  and AND2_0(G632,G62,G178);
  not NOT_0(G633,G164);
  not NOT_1(G634,G166);
  not NOT_2(G647,G167);
  not NOT_3(G659,G168);
  not NOT_4(G671,G169);
  nand NAND2_0(G684,G134,G1);
  not NOT_5(G685,G165);
  not NOT_6(G686,G632);
  and AND2_1(G687,G633,G11);
  and AND2_2(G688,G136,G154);
  and AND4_0(G689,G136,G155,G154,G153);
  not NOT_7(G690,G157);
  not NOT_8(G694,G158);
  not NOT_9(G706,G159);
  not NOT_10(G718,G158);
  not NOT_11(G730,G159);
  not NOT_12(G742,G64);
  not NOT_13(G746,G64);
  not NOT_14(G749,G66);
  not NOT_15(G752,G162);
  not NOT_16(G756,G160);
  not NOT_17(G768,G161);
  not NOT_18(G780,G160);
  not NOT_19(G792,G161);
  not NOT_20(G804,G102);
  not NOT_21(G813,G101);
  not NOT_22(G825,G101);
  not NOT_23(G836,G100);
  not NOT_24(G848,G100);
  not NOT_25(G860,G173);
  not NOT_26(G872,G172);
  not NOT_27(G884,G174);
  not NOT_28(G896,G175);
  not NOT_29(G908,G90);
  not NOT_30(G911,G90);
  not NOT_31(G914,G92);
  not NOT_32(G917,G92);
  not NOT_33(G920,G94);
  not NOT_34(G923,G94);
  not NOT_35(G926,G96);
  not NOT_36(G929,G96);
  not NOT_37(G932,G103);
  not NOT_38(G935,G103);
  not NOT_39(G938,G105);
  not NOT_40(G941,G105);
  not NOT_41(G944,G107);
  not NOT_42(G947,G107);
  not NOT_43(G950,G109);
  not NOT_44(G953,G109);
  not NOT_45(G956,G124);
  not NOT_46(G963,G124);
  not NOT_47(G970,G88);
  and AND2_3(G976,G11,G12);
  not NOT_48(G980,G1);
  not NOT_49(G983,G163);
  not NOT_50(G993,G113);
  not NOT_51(G996,G115);
  not NOT_52(G999,G117);
  not NOT_53(G1002,G117);
  not NOT_54(G1005,G119);
  not NOT_55(G1008,G119);
  not NOT_56(G1011,G121);
  not NOT_57(G1014,G121);
  not NOT_58(G1017,G126);
  not NOT_59(G1020,G126);
  not NOT_60(G1023,G128);
  not NOT_61(G1026,G128);
  not NOT_62(G1029,G103);
  not NOT_63(G1032,G103);
  not NOT_64(G1035,G105);
  not NOT_65(G1038,G105);
  not NOT_66(G1041,G107);
  not NOT_67(G1044,G107);
  not NOT_68(G1047,G109);
  not NOT_69(G1050,G109);
  not NOT_70(G1053,G123);
  not NOT_71(G1060,G123);
  not NOT_72(G1067,G152);
  and AND2_4(G1070,G12,G11);
  not NOT_73(G1075,G163);
  not NOT_74(G1081,G121);
  not NOT_75(G1084,G121);
  not NOT_76(G1087,G126);
  not NOT_77(G1090,G126);
  not NOT_78(G1093,G128);
  not NOT_79(G1096,G128);
  not NOT_80(G1099,G113);
  not NOT_81(G1102,G115);
  not NOT_82(G1105,G117);
  not NOT_83(G1108,G117);
  not NOT_84(G1111,G119);
  not NOT_85(G1114,G119);
  not NOT_86(G1117,G130);
  not NOT_87(G1120,G130);
  not NOT_88(G1123,G90);
  not NOT_89(G1126,G90);
  not NOT_90(G1129,G92);
  not NOT_91(G1132,G92);
  not NOT_92(G1135,G94);
  not NOT_93(G1138,G94);
  not NOT_94(G1141,G96);
  not NOT_95(G1144,G96);
  not NOT_96(G1147,G121);
  not NOT_97(G1150,G98);
  not NOT_98(G1162,G98);
  not NOT_99(G1172,G102);
  not NOT_100(G1184,G173);
  not NOT_101(G1196,G172);
  not NOT_102(G1208,G177);
  not NOT_103(G1214,G176);
  not NOT_104(G1218,G174);
  not NOT_105(G1230,G175);
  not NOT_106(G1242,G170);
  not NOT_107(G1245,G171);
  not NOT_108(G1248,G176);
  not NOT_109(G1256,G177);
  not NOT_110(G1264,G176);
  not NOT_111(G1272,G177);
  not NOT_112(G1280,G176);
  not NOT_113(G1287,G177);
  not NOT_114(G1294,G176);
  not NOT_115(G1301,G177);
  not NOT_116(G1308,G114);
  not NOT_117(G1311,G142);
  not NOT_118(G1314,G143);
  not NOT_119(G1317,G144);
  not NOT_120(G1320,G140);
  not NOT_121(G1323,G141);
  not NOT_122(G1326,G137);
  not NOT_123(G1329,G138);
  not NOT_124(G1332,G139);
  not NOT_125(G1335,G135);
  not NOT_126(G1338,G2);
  not NOT_127(G1341,G142);
  not NOT_128(G1344,G143);
  not NOT_129(G1347,G144);
  not NOT_130(G1350,G141);
  not NOT_131(G1353,G137);
  not NOT_132(G1356,G138);
  not NOT_133(G1359,G139);
  not NOT_134(G1362,G140);
  not NOT_135(G1365,G135);
  not NOT_136(G1368,G145);
  not NOT_137(G1371,G146);
  not NOT_138(G1374,G147);
  not NOT_139(G1377,G148);
  not NOT_140(G1380,G149);
  not NOT_141(G1383,G150);
  not NOT_142(G1386,G21);
  not NOT_143(G1389,G145);
  not NOT_144(G1392,G147);
  not NOT_145(G1395,G148);
  not NOT_146(G1398,G149);
  not NOT_147(G1401,G150);
  not NOT_148(G1404,G146);
  not NOT_149(G1407,G130);
  not NOT_150(G1410,G132);
  not NOT_151(G1413,G126);
  not NOT_152(G1416,G128);
  not NOT_153(G1419,G117);
  not NOT_154(G1422,G119);
  not NOT_155(G1425,G113);
  not NOT_156(G1428,G115);
  not NOT_157(G1431,G109);
  not NOT_158(G1434,G111);
  not NOT_159(G1437,G105);
  not NOT_160(G1440,G107);
  not NOT_161(G1443,G96);
  not NOT_162(G1446,G103);
  not NOT_163(G1449,G92);
  not NOT_164(G1452,G94);
  not NOT_165(G1455,G90);
  and AND2_5(G1458,G671,G148);
  or OR2_0(G1459,G634,G148);
  and AND3_0(G1460,G76,G694,G706);
  and AND3_1(G1461,G77,G694,G706);
  and AND3_2(G1462,G75,G694,G706);
  and AND3_3(G1463,G74,G694,G706);
  and AND3_4(G1464,G73,G694,G706);
  and AND3_5(G1465,G81,G718,G730);
  and AND3_6(G1466,G72,G718,G730);
  and AND3_7(G1467,G70,G718,G730);
  and AND3_8(G1468,G68,G718,G730);
  and AND3_9(G1469,G76,G756,G768);
  and AND3_10(G1470,G77,G756,G768);
  and AND3_11(G1471,G75,G756,G768);
  and AND3_12(G1472,G74,G756,G768);
  and AND3_13(G1473,G73,G756,G768);
  and AND3_14(G1474,G81,G780,G792);
  and AND3_15(G1475,G72,G780,G792);
  and AND3_16(G1476,G70,G780,G792);
  and AND3_17(G1477,G68,G780,G792);
  and AND3_18(G1478,G41,G1218,G1230);
  and AND3_19(G1479,G22,G860,G872);
  and AND3_20(G1480,G41,G1184,G1196);
  and AND3_21(G1481,G18,G1184,G1196);
  and AND3_22(G1482,G40,G1184,G1196);
  and AND3_23(G1483,G15,G1184,G1196);
  and AND3_24(G1484,G14,G1184,G1196);
  and AND3_25(G1485,G6,G860,G872);
  and AND3_26(G1486,G5,G860,G872);
  and AND3_27(G1487,G25,G860,G872);
  and AND3_28(G1488,G23,G860,G872);
  and AND3_29(G1489,G18,G1218,G1230);
  and AND3_30(G1490,G40,G1218,G1230);
  and AND3_31(G1491,G15,G1218,G1230);
  and AND3_32(G1492,G14,G1218,G1230);
  and AND3_33(G1493,G6,G884,G896);
  and AND3_34(G1494,G5,G884,G896);
  and AND3_35(G1495,G25,G884,G896);
  and AND3_36(G1496,G23,G884,G896);
  and AND3_37(G1497,G54,G1245,G170);
  and AND2_6(G1498,G1264,G1272);
  and AND3_38(G1499,G22,G884,G896);
  and AND2_7(G1500,G1248,G1256);
  not NOT_166(G1501,G1311);
  not NOT_167(G1502,G1314);
  not NOT_168(G1503,G1317);
  not NOT_169(G1504,G1320);
  not NOT_170(G1505,G1323);
  not NOT_171(G1506,G1326);
  not NOT_172(G1507,G1329);
  not NOT_173(G1508,G1332);
  not NOT_174(G1509,G1335);
  not NOT_175(G1510,G1338);
  not NOT_176(G1511,G1341);
  not NOT_177(G1512,G1344);
  not NOT_178(G1513,G1347);
  not NOT_179(G1514,G1350);
  not NOT_180(G1515,G1353);
  not NOT_181(G1516,G1356);
  not NOT_182(G1517,G1359);
  not NOT_183(G1518,G1362);
  not NOT_184(G1519,G1365);
  not NOT_185(G1520,G742);
  not NOT_186(G1526,G694);
  not NOT_187(G1537,G706);
  not NOT_188(G1548,G742);
  not NOT_189(G1554,G718);
  not NOT_190(G1565,G730);
  and AND3_39(G1576,G79,G718,G730);
  not NOT_191(G1577,G980);
  not NOT_192(G1582,G1368);
  not NOT_193(G1583,G1371);
  not NOT_194(G1584,G1374);
  not NOT_195(G1585,G1377);
  not NOT_196(G1586,G1380);
  not NOT_197(G1587,G1383);
  not NOT_198(G1588,G1386);
  not NOT_199(G1589,G1389);
  not NOT_200(G1590,G1392);
  not NOT_201(G1591,G1395);
  not NOT_202(G1592,G1398);
  not NOT_203(G1593,G1401);
  not NOT_204(G1594,G1404);
  not NOT_205(G1595,G746);
  not NOT_206(G1601,G756);
  not NOT_207(G1612,G768);
  not NOT_208(G1623,G746);
  not NOT_209(G1629,G780);
  not NOT_210(G1640,G792);
  and AND3_40(G1651,G79,G780,G792);
  not NOT_211(G1652,G860);
  not NOT_212(G1663,G872);
  not NOT_213(G1674,G884);
  not NOT_214(G1685,G896);
  not NOT_215(G1696,G908);
  not NOT_216(G1697,G911);
  not NOT_217(G1698,G914);
  not NOT_218(G1699,G917);
  not NOT_219(G1700,G920);
  not NOT_220(G1701,G923);
  not NOT_221(G1702,G926);
  not NOT_222(G1703,G929);
  and AND3_41(G1704,G671,G143,G911);
  and AND3_42(G1705,G671,G144,G917);
  and AND3_43(G1706,G671,G140,G923);
  and AND3_44(G1707,G671,G141,G929);
  and AND2_8(G1708,G634,G908);
  and AND2_9(G1709,G634,G914);
  and AND2_10(G1710,G634,G920);
  and AND2_11(G1711,G634,G926);
  not NOT_223(G1712,G932);
  not NOT_224(G1713,G935);
  not NOT_225(G1714,G938);
  not NOT_226(G1715,G941);
  not NOT_227(G1716,G944);
  not NOT_228(G1717,G947);
  not NOT_229(G1718,G950);
  not NOT_230(G1719,G953);
  and AND3_45(G1720,G671,G137,G935);
  and AND3_46(G1721,G671,G138,G941);
  and AND3_47(G1722,G671,G139,G947);
  and AND3_48(G1723,G671,G135,G953);
  and AND2_12(G1724,G634,G932);
  and AND2_13(G1725,G634,G938);
  and AND2_14(G1726,G634,G944);
  and AND2_15(G1727,G634,G950);
  not NOT_231(G1728,G956);
  not NOT_232(G1734,G963);
  and AND2_16(G1740,G112,G956);
  and AND2_17(G1741,G110,G956);
  and AND2_18(G1742,G108,G956);
  and AND2_19(G1743,G106,G956);
  and AND2_20(G1744,G104,G956);
  and AND2_21(G1745,G97,G963);
  and AND2_22(G1746,G95,G963);
  and AND2_23(G1747,G93,G963);
  and AND2_24(G1748,G91,G963);
  and AND2_25(G1749,G89,G963);
  not NOT_233(G1750,G749);
  not NOT_234(G1755,G983);
  not NOT_235(G1764,G976);
  not NOT_236(G1774,G993);
  not NOT_237(G1775,G996);
  not NOT_238(G1776,G999);
  not NOT_239(G1777,G1002);
  not NOT_240(G1778,G1005);
  not NOT_241(G1779,G1008);
  and AND2_26(G1780,G836,G996);
  and AND3_49(G1781,G836,G145,G1002);
  and AND3_50(G1782,G836,G146,G1008);
  and AND2_27(G1783,G1150,G993);
  and AND2_28(G1784,G1150,G999);
  and AND2_29(G1785,G1150,G1005);
  not NOT_242(G1786,G1011);
  not NOT_243(G1787,G1014);
  not NOT_244(G1788,G1017);
  not NOT_245(G1789,G1020);
  not NOT_246(G1790,G1023);
  not NOT_247(G1791,G1026);
  and AND3_51(G1792,G671,G147,G1014);
  not NOT_248(G1793,G1458);
  and AND3_52(G1794,G671,G149,G1020);
  and AND3_53(G1795,G671,G150,G1026);
  and AND2_30(G1796,G634,G1011);
  and AND2_31(G1797,G634,G1017);
  and AND2_32(G1798,G634,G1023);
  not NOT_249(G1799,G1029);
  not NOT_250(G1800,G1032);
  not NOT_251(G1801,G1035);
  not NOT_252(G1802,G1038);
  not NOT_253(G1803,G1041);
  not NOT_254(G1804,G1044);
  not NOT_255(G1805,G1047);
  not NOT_256(G1806,G1050);
  and AND3_54(G1807,G836,G137,G1032);
  and AND3_55(G1808,G836,G138,G1038);
  and AND3_56(G1809,G836,G139,G1044);
  and AND3_57(G1810,G836,G135,G1050);
  and AND2_33(G1811,G1150,G1029);
  and AND2_34(G1812,G1150,G1035);
  and AND2_35(G1813,G1150,G1041);
  and AND2_36(G1814,G1150,G1047);
  not NOT_257(G1815,G1053);
  not NOT_258(G1821,G1060);
  and AND2_37(G1827,G133,G1053);
  and AND2_38(G1828,G131,G1053);
  and AND2_39(G1829,G129,G1053);
  and AND2_40(G1830,G127,G1053);
  and AND2_41(G1831,G125,G1053);
  and AND2_42(G1832,G122,G1060);
  and AND2_43(G1833,G120,G1060);
  and AND2_44(G1834,G118,G1060);
  and AND2_45(G1835,G116,G1060);
  and AND2_46(G1836,G114,G1060);
  not NOT_259(G1837,G1075);
  and AND2_47(G1842,G32,G1075);
  and AND2_48(G1843,G33,G1075);
  and AND2_49(G1844,G35,G1075);
  and AND2_50(G1845,G35,G1075);
  not NOT_260(G1846,G1081);
  not NOT_261(G1847,G1084);
  not NOT_262(G1848,G1087);
  not NOT_263(G1849,G1090);
  not NOT_264(G1850,G1093);
  not NOT_265(G1851,G1096);
  and AND3_58(G1852,G848,G147,G1084);
  and AND2_51(G1853,G848,G148);
  and AND3_59(G1854,G848,G149,G1090);
  and AND3_60(G1855,G848,G150,G1096);
  and AND2_52(G1856,G1162,G1081);
  or OR2_1(G1857,G1162,G148);
  and AND2_53(G1858,G1162,G1087);
  and AND2_54(G1859,G1162,G1093);
  not NOT_266(G1860,G1099);
  not NOT_267(G1861,G1102);
  not NOT_268(G1862,G1105);
  not NOT_269(G1863,G1108);
  not NOT_270(G1864,G1111);
  not NOT_271(G1865,G1114);
  and AND2_55(G1866,G848,G1102);
  and AND3_61(G1867,G848,G145,G1108);
  and AND3_62(G1868,G848,G146,G1114);
  and AND2_56(G1869,G1162,G1099);
  and AND2_57(G1870,G1162,G1105);
  and AND2_58(G1871,G1162,G1111);
  not NOT_272(G1872,G1117);
  not NOT_273(G1873,G970);
  not NOT_274(G1876,G970);
  not NOT_275(G1879,G1120);
  not NOT_276(G1880,G970);
  not NOT_277(G1883,G970);
  and AND2_59(G1886,G848,G1117);
  and AND2_60(G1887,G848,G1120);
  not NOT_278(G1888,G1123);
  not NOT_279(G1889,G1126);
  not NOT_280(G1890,G1129);
  not NOT_281(G1891,G1132);
  not NOT_282(G1892,G1135);
  not NOT_283(G1893,G1138);
  not NOT_284(G1894,G1141);
  not NOT_285(G1895,G1144);
  and AND3_63(G1896,G836,G143,G1126);
  and AND3_64(G1897,G836,G144,G1132);
  and AND3_65(G1898,G836,G140,G1138);
  and AND3_66(G1899,G836,G141,G1144);
  and AND2_61(G1900,G1150,G1123);
  and AND2_62(G1901,G1150,G1129);
  and AND2_63(G1902,G1150,G1135);
  and AND2_64(G1903,G1150,G1141);
  not NOT_286(G1904,G1407);
  not NOT_287(G1905,G1410);
  not NOT_288(G1906,G1413);
  not NOT_289(G1907,G1416);
  not NOT_290(G1908,G1147);
  not NOT_291(G1911,G1147);
  not NOT_292(G1914,G1184);
  not NOT_293(G1925,G1196);
  not NOT_294(G1936,G1208);
  not NOT_295(G1941,G1214);
  and AND2_65(G1944,G38,G1208);
  and AND2_66(G1945,G37,G1208);
  and AND2_67(G1946,G38,G1208);
  and AND2_68(G1947,G37,G1208);
  not NOT_296(G1948,G1218);
  not NOT_297(G1959,G1230);
  not NOT_298(G1970,G1248);
  not NOT_299(G1981,G1256);
  not NOT_300(G1992,G1264);
  not NOT_301(G2003,G1272);
  not NOT_302(G2014,G1431);
  not NOT_303(G2015,G1434);
  not NOT_304(G2016,G1437);
  not NOT_305(G2017,G1440);
  not NOT_306(G2018,G1443);
  not NOT_307(G2019,G1446);
  not NOT_308(G2020,G1280);
  not NOT_309(G2031,G1287);
  not NOT_310(G2042,G1294);
  not NOT_311(G2053,G1301);
  not NOT_312(G2064,G1308);
  not NOT_313(G2067,G1419);
  not NOT_314(G2068,G1422);
  not NOT_315(G2069,G1425);
  not NOT_316(G2070,G1428);
  not NOT_317(G2071,G1449);
  not NOT_318(G2072,G1452);
  not NOT_319(G2073,G970);
  not NOT_320(G2076,G1455);
  and AND3_67(G2077,G143,G659,G1697);
  and AND3_68(G2078,G144,G659,G1699);
  and AND3_69(G2079,G140,G659,G1701);
  and AND3_70(G2080,G141,G659,G1703);
  and AND2_69(G2081,G647,G1696);
  and AND2_70(G2082,G647,G1698);
  and AND2_71(G2083,G647,G1700);
  and AND2_72(G2084,G647,G1702);
  and AND3_71(G2085,G137,G659,G1713);
  and AND3_72(G2086,G138,G659,G1715);
  and AND3_73(G2087,G139,G659,G1717);
  and AND3_74(G2088,G135,G659,G1719);
  and AND2_73(G2089,G647,G1712);
  and AND2_74(G2090,G647,G1714);
  and AND2_75(G2091,G647,G1716);
  and AND2_76(G2092,G647,G1718);
  and AND2_77(G2093,G813,G1775);
  and AND3_75(G2094,G145,G813,G1777);
  and AND3_76(G2095,G146,G813,G1779);
  and AND2_78(G2096,G1172,G1774);
  and AND2_79(G2097,G1172,G1776);
  and AND2_80(G2098,G1172,G1778);
  and AND3_77(G2099,G147,G659,G1787);
  and AND3_78(G2100,G149,G659,G1789);
  and AND3_79(G2101,G150,G659,G1791);
  and AND2_81(G2102,G647,G1786);
  and AND2_82(G2103,G647,G1788);
  and AND2_83(G2104,G647,G1790);
  and AND2_84(G2105,G1793,G1459);
  and AND3_80(G2108,G137,G813,G1800);
  and AND3_81(G2109,G138,G813,G1802);
  and AND3_82(G2110,G139,G813,G1804);
  and AND3_83(G2111,G135,G813,G1806);
  and AND2_85(G2112,G1172,G1799);
  and AND2_86(G2113,G1172,G1801);
  and AND2_87(G2114,G1172,G1803);
  and AND2_88(G2115,G1172,G1805);
  and AND3_84(G2116,G147,G825,G1847);
  not NOT_321(G2117,G1853);
  and AND3_85(G2118,G149,G825,G1849);
  and AND3_86(G2119,G150,G825,G1851);
  and AND2_89(G2120,G804,G1846);
  and AND2_90(G2121,G804,G1848);
  and AND2_91(G2122,G804,G1850);
  and AND2_92(G2123,G825,G1861);
  and AND3_87(G2124,G145,G825,G1863);
  and AND3_88(G2125,G146,G825,G1865);
  and AND2_93(G2126,G804,G1860);
  and AND2_94(G2127,G804,G1862);
  and AND2_95(G2128,G804,G1864);
  and AND2_96(G2129,G825,G1872);
  and AND2_97(G2130,G825,G1879);
  and AND3_89(G2131,G143,G813,G1889);
  and AND3_90(G2132,G144,G813,G1891);
  and AND3_91(G2133,G140,G813,G1893);
  and AND3_92(G2134,G141,G813,G1895);
  and AND2_98(G2135,G1172,G1888);
  and AND2_99(G2136,G1172,G1890);
  and AND2_100(G2137,G1172,G1892);
  and AND2_101(G2138,G1172,G1894);
  nand NAND2_1(G2139,G1410,G1904);
  nand NAND2_2(G2140,G1407,G1905);
  nand NAND2_3(G2141,G1416,G1906);
  nand NAND2_4(G2142,G1413,G1907);
  nand NAND2_5(G2143,G1434,G2014);
  nand NAND2_6(G2144,G1431,G2015);
  nand NAND2_7(G2145,G1440,G2016);
  nand NAND2_8(G2146,G1437,G2017);
  nand NAND2_9(G2147,G1446,G2018);
  nand NAND2_10(G2148,G1443,G2019);
  nand NAND2_11(G2149,G1422,G2067);
  nand NAND2_12(G2150,G1419,G2068);
  nand NAND2_13(G2151,G1428,G2069);
  nand NAND2_14(G2152,G1425,G2070);
  nand NAND2_15(G2153,G1452,G2071);
  nand NAND2_16(G2154,G1449,G2072);
  and AND2_102(G2155,G1755,G1764);
  and AND2_103(G2156,G983,G1764);
  and AND3_93(G2157,G86,G1526,G706);
  and AND3_94(G2158,G87,G1526,G706);
  and AND3_95(G2159,G85,G1526,G706);
  and AND3_96(G2160,G84,G1526,G706);
  and AND3_97(G2161,G83,G1526,G706);
  and AND3_98(G2162,G80,G1554,G730);
  and AND3_99(G2163,G82,G1554,G730);
  and AND3_100(G2164,G71,G1554,G730);
  and AND3_101(G2165,G69,G1554,G730);
  and AND2_104(G2166,G1755,G1764);
  and AND2_105(G2167,G983,G1764);
  and AND3_102(G2168,G86,G1601,G768);
  and AND3_103(G2169,G87,G1601,G768);
  and AND3_104(G2170,G85,G1601,G768);
  and AND3_105(G2171,G84,G1601,G768);
  and AND3_106(G2172,G83,G1601,G768);
  and AND3_107(G2173,G80,G1629,G792);
  and AND3_108(G2174,G82,G1629,G792);
  and AND3_109(G2175,G71,G1629,G792);
  and AND3_110(G2176,G69,G1629,G792);
  and AND2_106(G2177,G1755,G1764);
  and AND2_107(G2178,G983,G1764);
  and AND3_111(G2179,G42,G1948,G1230);
  and AND2_108(G2180,G1755,G1764);
  and AND2_109(G2181,G983,G1764);
  and AND3_112(G2182,G3,G1652,G872);
  and AND3_113(G2183,G42,G1914,G1196);
  and AND3_114(G2184,G17,G1914,G1196);
  and AND3_115(G2185,G39,G1914,G1196);
  and AND3_116(G2186,G36,G1914,G1196);
  and AND3_117(G2187,G16,G1914,G1196);
  and AND3_118(G2188,G27,G1652,G872);
  and AND3_119(G2189,G26,G1652,G872);
  and AND3_120(G2190,G24,G1652,G872);
  and AND3_121(G2191,G4,G1652,G872);
  and AND3_122(G2192,G17,G1948,G1230);
  and AND3_123(G2193,G39,G1948,G1230);
  and AND3_124(G2194,G36,G1948,G1230);
  and AND3_125(G2195,G16,G1948,G1230);
  and AND3_126(G2196,G27,G1674,G896);
  and AND3_127(G2197,G26,G1674,G896);
  and AND3_128(G2198,G24,G1674,G896);
  and AND3_129(G2199,G4,G1674,G896);
  and AND3_130(G2200,G51,G1992,G1272);
  and AND3_131(G2201,G3,G1674,G896);
  and AND3_132(G2202,G49,G1970,G1256);
  and AND3_133(G2203,G78,G1554,G730);
  and AND3_134(G2204,G78,G1629,G792);
  or OR2_2(G2205,G1704,G2077);
  or OR2_3(G2206,G1705,G2078);
  or OR2_4(G2207,G1706,G2079);
  or OR2_5(G2208,G1707,G2080);
  or OR3_0(G2209,G1708,G2081,G143);
  or OR3_1(G2210,G1709,G2082,G144);
  or OR3_2(G2211,G1710,G2083,G140);
  or OR3_3(G2212,G1711,G2084,G141);
  or OR2_6(G2213,G1720,G2085);
  or OR2_7(G2214,G1721,G2086);
  or OR2_8(G2215,G1722,G2087);
  or OR2_9(G2216,G1723,G2088);
  or OR3_4(G2217,G1724,G2089,G137);
  or OR3_5(G2218,G1725,G2090,G138);
  or OR3_6(G2219,G1726,G2091,G139);
  or OR3_7(G2220,G1727,G2092,G135);
  and AND2_110(G2221,G111,G1728);
  and AND2_111(G2222,G109,G1728);
  and AND2_112(G2223,G107,G1728);
  and AND2_113(G2224,G105,G1728);
  and AND2_114(G2225,G103,G1728);
  and AND2_115(G2226,G96,G1734);
  and AND2_116(G2227,G94,G1734);
  and AND2_117(G2228,G92,G1734);
  and AND2_118(G2229,G90,G1734);
  and AND2_119(G2230,G88,G1734);
  not NOT_322(G2231,G1764);
  or OR2_10(G2240,G1780,G2093);
  or OR2_11(G2241,G1781,G2094);
  or OR2_12(G2242,G1782,G2095);
  or OR3_8(G2243,G1784,G2097,G145);
  or OR3_9(G2244,G1785,G2098,G146);
  or OR2_13(G2245,G1783,G2096);
  or OR2_14(G2248,G1792,G2099);
  or OR2_15(G2249,G1794,G2100);
  or OR2_16(G2250,G1795,G2101);
  or OR3_10(G2251,G1796,G2102,G147);
  or OR3_11(G2252,G1797,G2103,G149);
  or OR3_12(G2253,G1798,G2104,G150);
  or OR2_17(G2254,G1807,G2108);
  or OR2_18(G2255,G1808,G2109);
  or OR2_19(G2256,G1809,G2110);
  or OR2_20(G2257,G1810,G2111);
  or OR3_13(G2258,G1811,G2112,G137);
  or OR3_14(G2259,G1812,G2113,G138);
  or OR3_15(G2260,G1813,G2114,G139);
  or OR3_16(G2261,G1814,G2115,G135);
  and AND2_120(G2262,G132,G1815);
  and AND2_121(G2263,G130,G1815);
  and AND2_122(G2264,G128,G1815);
  and AND2_123(G2265,G126,G1815);
  and AND2_124(G2266,G121,G1821);
  and AND2_125(G2267,G119,G1821);
  and AND2_126(G2268,G117,G1821);
  and AND2_127(G2269,G115,G1821);
  and AND2_128(G2270,G113,G1821);
  or OR2_21(G2271,G1815,G1831);
  and AND2_129(G2277,G32,G1837);
  and AND2_130(G2278,G34,G1837);
  and AND2_131(G2279,G13,G1837);
  and AND2_132(G2280,G13,G1837);
  or OR2_22(G2281,G1852,G2116);
  or OR2_23(G2282,G1854,G2118);
  or OR2_24(G2283,G1855,G2119);
  or OR3_17(G2284,G1856,G2120,G147);
  or OR3_18(G2285,G1858,G2121,G149);
  or OR3_19(G2286,G1859,G2122,G150);
  or OR2_25(G2287,G1866,G2123);
  or OR2_26(G2288,G1867,G2124);
  or OR2_27(G2289,G1868,G2125);
  or OR3_20(G2290,G1870,G2127,G145);
  or OR3_21(G2291,G1871,G2128,G146);
  not NOT_323(G2292,G1873);
  not NOT_324(G2293,G1876);
  not NOT_325(G2294,G1880);
  not NOT_326(G2295,G1883);
  or OR2_28(G2296,G1886,G2129);
  and AND3_135(G2297,G848,G142,G1876);
  or OR2_29(G2298,G1887,G2130);
  and AND3_136(G2299,G848,G142,G1883);
  and AND2_133(G2300,G1162,G1873);
  and AND2_134(G2301,G1162,G1880);
  or OR2_30(G2302,G1896,G2131);
  or OR2_31(G2303,G1897,G2132);
  or OR2_32(G2304,G1898,G2133);
  or OR2_33(G2305,G1899,G2134);
  or OR3_22(G2306,G1900,G2135,G143);
  or OR3_23(G2307,G1901,G2136,G144);
  or OR3_24(G2308,G1902,G2137,G140);
  or OR3_25(G2309,G1903,G2138,G141);
  nand NAND2_17(G2310,G2139,G2140);
  nand NAND2_18(G2314,G2141,G2142);
  not NOT_327(G2318,G1908);
  not NOT_328(G2319,G1911);
  and AND3_137(G2320,G48,G1970,G1256);
  and AND3_138(G2321,G55,G1970,G1256);
  and AND3_139(G2322,G56,G1970,G1256);
  and AND3_140(G2323,G57,G1970,G1256);
  and AND3_141(G2324,G60,G1992,G1272);
  and AND3_142(G2325,G58,G1992,G1272);
  and AND3_143(G2326,G50,G1992,G1272);
  and AND3_144(G2327,G59,G1992,G1272);
  nand NAND2_19(G2328,G2143,G2144);
  nand NAND2_20(G2332,G2145,G2146);
  nand NAND2_21(G2336,G2147,G2148);
  and AND3_145(G2339,G53,G2020,G1287);
  and AND3_146(G2340,G44,G2020,G1287);
  and AND3_147(G2341,G20,G2020,G1287);
  and AND3_148(G2342,G45,G2020,G1287);
  and AND3_149(G2343,G46,G2020,G1287);
  and AND3_150(G2344,G19,G2042,G1301);
  and AND3_151(G2345,G43,G2042,G1301);
  and AND3_152(G2346,G47,G2042,G1301);
  and AND3_153(G2347,G52,G2042,G1301);
  and AND3_154(G2348,G54,G2042,G1301);
  nand NAND2_22(G2349,G2151,G2152);
  nand NAND2_23(G2352,G2149,G2150);
  and AND2_135(G2355,G2117,G1857);
  or OR2_34(G2358,G1869,G2126);
  not NOT_329(G2361,G2073);
  nand NAND2_24(G2362,G2073,G2076);
  nand NAND2_25(G2363,G2153,G2154);
  not NOT_330(G2366,G2105);
  or OR2_35(G2367,G2278,G1843);
  or OR2_36(G2368,G2279,G1844);
  or OR2_37(G2369,G2280,G1845);
  or OR2_38(G2370,G2277,G1842);
  not NOT_331(G2371,G2205);
  not NOT_332(G2372,G2206);
  not NOT_333(G2373,G2207);
  not NOT_334(G2374,G2208);
  not NOT_335(G2375,G2213);
  not NOT_336(G2376,G2214);
  not NOT_337(G2377,G2215);
  not NOT_338(G2378,G2216);
  or OR2_39(G2379,G2222,G1741);
  or OR2_40(G2386,G2223,G1742);
  or OR2_41(G2392,G2224,G1743);
  or OR2_42(G2398,G2225,G1744);
  or OR2_43(G2404,G2226,G1745);
  or OR2_44(G2410,G2227,G1746);
  or OR2_45(G2418,G2228,G1747);
  or OR2_46(G2424,G2229,G1748);
  or OR2_47(G2430,G2230,G1749);
  not NOT_339(G2436,G2241);
  not NOT_340(G2437,G2242);
  not NOT_341(G2438,G2240);
  not NOT_342(G2441,G2248);
  not NOT_343(G2442,G2249);
  not NOT_344(G2443,G2250);
  not NOT_345(G2444,G2254);
  not NOT_346(G2445,G2255);
  not NOT_347(G2446,G2256);
  not NOT_348(G2447,G2257);
  or OR2_48(G2448,G2263,G1828);
  or OR2_49(G2454,G2264,G1829);
  or OR2_50(G2460,G2265,G1830);
  or OR2_51(G2466,G2266,G1832);
  or OR2_52(G2472,G2267,G1833);
  or OR2_53(G2480,G2268,G1834);
  or OR2_54(G2486,G2269,G1835);
  or OR2_55(G2492,G2270,G1836);
  not NOT_349(G2499,G2281);
  not NOT_350(G2500,G2282);
  not NOT_351(G2501,G2283);
  not NOT_352(G2502,G2288);
  not NOT_353(G2503,G2289);
  and AND3_155(G2504,G142,G825,G2293);
  and AND3_156(G2505,G142,G825,G2295);
  and AND2_136(G2506,G804,G2292);
  and AND2_137(G2507,G804,G2294);
  not NOT_354(G2508,G2296);
  not NOT_355(G2511,G2298);
  not NOT_356(G2512,G2302);
  not NOT_357(G2513,G2303);
  not NOT_358(G2514,G2304);
  not NOT_359(G2515,G2305);
  and AND3_157(G2516,G2105,G1992,G2003);
  or OR2_56(G2517,G2262,G1827);
  or OR2_57(G2520,G2221,G1740);
  not NOT_360(G2523,G2287);
  nand NAND2_26(G2526,G1455,G2361);
  not NOT_361(G2527,G2245);
  and AND2_138(G2528,G2367,G1070);
  and AND3_158(G2529,G8,G1755,G2231);
  and AND3_159(G2530,G9,G983,G2231);
  and AND3_160(G2531,G10,G1755,G2231);
  and AND3_161(G2532,G30,G983,G2231);
  and AND2_139(G2533,G2368,G1070);
  and AND3_162(G2534,G28,G1755,G2231);
  and AND3_163(G2535,G7,G983,G2231);
  and AND3_164(G2536,G31,G1755,G2231);
  and AND3_165(G2537,G29,G983,G2231);
  and AND2_140(G2538,G2369,G1070);
  and AND2_141(G2539,G2370,G1070);
  and AND2_142(G2540,G2271,G148);
  and AND2_143(G2543,G148,G2271);
  and AND2_144(G2547,G2371,G2209);
  and AND2_145(G2550,G2372,G2210);
  and AND2_146(G2553,G2373,G2211);
  and AND2_147(G2556,G2374,G2212);
  and AND2_148(G2559,G2375,G2217);
  and AND2_149(G2562,G2376,G2218);
  and AND2_150(G2565,G2377,G2219);
  and AND2_151(G2568,G2378,G2220);
  and AND2_152(G2571,G2436,G2243);
  and AND2_153(G2574,G2437,G2244);
  not NOT_362(G2577,G2245);
  and AND2_154(G2580,G2441,G2251);
  and AND2_155(G2583,G2442,G2252);
  and AND2_156(G2586,G2443,G2253);
  or OR2_58(G2589,G2297,G2504);
  or OR2_59(G2590,G2299,G2505);
  or OR3_26(G2591,G2300,G2506,G142);
  or OR3_27(G2592,G2301,G2507,G142);
  not NOT_363(G2593,G2310);
  not NOT_364(G2596,G2314);
  and AND3_166(G2599,G2314,G2310,G1908);
  and AND3_167(G2600,G2511,G1992,G2003);
  and AND2_157(G2601,G2447,G2261);
  not NOT_365(G2602,G2355);
  not NOT_366(G2603,G2328);
  not NOT_367(G2606,G2332);
  not NOT_368(G2609,G2336);
  not NOT_369(G2612,G2336);
  not NOT_370(G2615,G2271);
  not NOT_371(G2618,G2271);
  not NOT_372(G2621,G2271);
  not NOT_373(G2624,G2349);
  not NOT_374(G2625,G2352);
  and AND2_158(G2626,G2445,G2259);
  and AND2_159(G2629,G2446,G2260);
  and AND2_160(G2632,G2515,G2309);
  and AND2_161(G2635,G2444,G2258);
  and AND2_162(G2638,G2513,G2307);
  and AND2_163(G2641,G2514,G2308);
  and AND2_164(G2644,G2512,G2306);
  and AND2_165(G2647,G2500,G2285);
  and AND2_166(G2650,G2501,G2286);
  and AND2_167(G2653,G2499,G2284);
  and AND2_168(G2656,G2502,G2290);
  and AND2_169(G2659,G2503,G2291);
  not NOT_375(G2662,G2358);
  nand NAND2_27(G2663,G2526,G2362);
  not NOT_376(G2666,G2363);
  and AND2_170(G2667,G142,G2430);
  not NOT_377(G2668,G2438);
  not NOT_378(G2669,G2508);
  and AND2_171(G2670,G2430,G142);
  or OR4_0(G2671,G2529,G2530,G2155,G2156);
  or OR4_1(G2672,G2531,G2532,G2166,G2167);
  or OR4_2(G2673,G2534,G2535,G2177,G2178);
  or OR4_3(G2674,G2536,G2537,G2180,G2181);
  and AND2_172(G2675,G2424,G143);
  and AND2_173(G2679,G2418,G144);
  and AND2_174(G2685,G140,G2410);
  and AND2_175(G2692,G2404,G141);
  and AND2_176(G2693,G2398,G137);
  and AND2_177(G2696,G2392,G138);
  and AND2_178(G2700,G2386,G139);
  and AND2_179(G2705,G2379,G135);
  and AND2_180(G2711,G143,G2424);
  and AND2_181(G2715,G144,G2418);
  and AND2_182(G2720,G140,G2410);
  and AND2_183(G2726,G141,G2404);
  and AND2_184(G2727,G137,G2398);
  and AND2_185(G2731,G138,G2392);
  and AND2_186(G2737,G139,G2386);
  and AND2_187(G2744,G135,G2379);
  not NOT_379(G2752,G2492);
  not NOT_380(G2759,G2486);
  not NOT_381(G2770,G2486);
  and AND2_188(G2774,G2480,G145);
  and AND2_189(G2780,G146,G2472);
  and AND2_190(G2787,G2466,G147);
  and AND2_191(G2788,G2460,G149);
  and AND2_192(G2792,G2454,G150);
  not NOT_382(G2797,G2448);
  not NOT_383(G2804,G2448);
  not NOT_384(G2810,G2492);
  not NOT_385(G2817,G2486);
  not NOT_386(G2828,G2486);
  and AND2_193(G2832,G145,G2480);
  and AND2_194(G2837,G146,G2472);
  and AND2_195(G2843,G147,G2466);
  and AND2_196(G2844,G149,G2460);
  and AND2_197(G2850,G150,G2454);
  not NOT_387(G2857,G2448);
  not NOT_388(G2865,G2448);
  not NOT_389(G2872,G2492);
  not NOT_390(G2875,G2589);
  not NOT_391(G2876,G2590);
  not NOT_392(G2877,G2517);
  not NOT_393(G2878,G2520);
  not NOT_394(G2879,G2601);
  not NOT_395(G2883,G2508);
  and AND3_168(G2887,G2438,G2042,G2053);
  not NOT_396(G2888,G2430);
  not NOT_397(G2891,G2424);
  not NOT_398(G2894,G2418);
  not NOT_399(G2897,G2410);
  not NOT_400(G2900,G2404);
  not NOT_401(G2903,G2398);
  not NOT_402(G2906,G2392);
  not NOT_403(G2909,G2386);
  not NOT_404(G2912,G2379);
  nor NOR2_0(G2915,G140,G2410);
  not NOT_405(G2918,G2430);
  not NOT_406(G2921,G2424);
  not NOT_407(G2924,G2418);
  not NOT_408(G2927,G2404);
  not NOT_409(G2930,G2398);
  not NOT_410(G2933,G2392);
  not NOT_411(G2936,G2386);
  not NOT_412(G2939,G2410);
  not NOT_413(G2942,G2379);
  nor NOR2_1(G2945,G140,G2410);
  nor NOR2_2(G2948,G135,G2379);
  not NOT_414(G2951,G2480);
  not NOT_415(G2954,G2472);
  not NOT_416(G2957,G2466);
  not NOT_417(G2960,G2460);
  not NOT_418(G2963,G2454);
  nor NOR2_3(G2966,G146,G2472);
  not NOT_419(G2969,G2480);
  not NOT_420(G2972,G2466);
  not NOT_421(G2975,G2460);
  not NOT_422(G2978,G2454);
  not NOT_423(G2981,G2472);
  nor NOR2_4(G2984,G146,G2472);
  not NOT_424(G2987,G2454);
  not NOT_425(G2990,G2460);
  not NOT_426(G2993,G2448);
  not NOT_427(G2996,G2466);
  not NOT_428(G2999,G2480);
  not NOT_429(G3002,G2472);
  not NOT_430(G3005,G2492);
  not NOT_431(G3008,G2486);
  not NOT_432(G3011,G2410);
  not NOT_433(G3014,G2404);
  not NOT_434(G3017,G2424);
  not NOT_435(G3020,G2418);
  not NOT_436(G3023,G2430);
  not NOT_437(G3026,G2386);
  not NOT_438(G3029,G2379);
  not NOT_439(G3032,G2398);
  not NOT_440(G3035,G2392);
  nand NAND2_28(G3038,G2352,G2624);
  nand NAND2_29(G3039,G2349,G2625);
  not NOT_441(G3040,G2523);
  nand NAND2_30(G3041,G2523,G2662);
  not NOT_442(G3042,G2574);
  not NOT_443(G3043,G2571);
  not NOT_444(G3044,G2586);
  not NOT_445(G3045,G2583);
  not NOT_446(G3046,G2580);
  not NOT_447(G3047,G2556);
  not NOT_448(G3048,G2553);
  not NOT_449(G3049,G2550);
  not NOT_450(G3050,G2547);
  not NOT_451(G3051,G2568);
  not NOT_452(G3052,G2565);
  not NOT_453(G3053,G2562);
  not NOT_454(G3054,G2559);
  and AND3_169(G3055,G2577,G1245,G1242);
  not NOT_455(G3056,G2615);
  nand NAND2_31(G3057,G2615,G1585);
  nand NAND2_32(G3058,G2618,G1591);
  not NOT_456(G3059,G2618);
  and AND2_198(G3060,G2875,G2591);
  and AND2_199(G3063,G2876,G2592);
  not NOT_457(G3064,G2621);
  and AND3_170(G3065,G2593,G2314,G2318);
  and AND3_171(G3066,G2310,G2596,G2319);
  and AND3_172(G3067,G2596,G2593,G1911);
  and AND3_173(G3068,G2568,G1970,G1981);
  and AND3_174(G3069,G2565,G1970,G1981);
  and AND3_175(G3070,G2562,G1970,G1981);
  and AND3_176(G3071,G2559,G1970,G1981);
  and AND3_177(G3072,G2586,G1992,G2003);
  and AND3_178(G3073,G2583,G1992,G2003);
  not NOT_458(G3074,G2626);
  not NOT_459(G3075,G2629);
  not NOT_460(G3076,G2632);
  not NOT_461(G3077,G2635);
  not NOT_462(G3078,G2647);
  not NOT_463(G3079,G2650);
  not NOT_464(G3080,G2653);
  nand NAND2_33(G3081,G2653,G2602);
  not NOT_465(G3082,G2609);
  not NOT_466(G3083,G2612);
  and AND3_179(G3084,G2332,G2328,G2609);
  and AND3_180(G3085,G2606,G2603,G2612);
  and AND3_181(G3086,G2556,G2020,G2031);
  and AND3_182(G3087,G2553,G2020,G2031);
  and AND3_183(G3088,G2550,G2020,G2031);
  and AND3_184(G3089,G2547,G2020,G2031);
  and AND3_185(G3090,G2580,G2042,G2053);
  and AND3_186(G3091,G2574,G2042,G2053);
  and AND3_187(G3092,G2571,G2042,G2053);
  and AND3_188(G3093,G2577,G2042,G2053);
  nand NAND2_34(G3094,G3038,G3039);
  not NOT_467(G3097,G2638);
  not NOT_468(G3098,G2641);
  not NOT_469(G3099,G2644);
  not NOT_470(G3100,G2656);
  not NOT_471(G3101,G2659);
  nand NAND2_35(G3102,G2358,G3040);
  not NOT_472(G3103,G2663);
  nand NAND2_36(G3104,G2663,G2666);
  and AND4_1(G3105,G3042,G3043,G2668,G2527);
  and AND4_2(G3106,G3044,G3045,G2366,G3046);
  and AND4_3(G3107,G3047,G3048,G3049,G3050);
  and AND4_4(G3108,G3051,G3052,G3053,G3054);
  and AND2_200(G3109,G2752,G2770);
  and AND3_189(G3110,G2759,G2752,G2774);
  and AND2_201(G3111,G2810,G2828);
  and AND3_190(G3112,G2817,G2810,G2832);
  not NOT_473(G3113,G2888);
  nand NAND2_37(G3114,G2888,G1501);
  not NOT_474(G3115,G2891);
  nand NAND2_38(G3116,G2891,G1502);
  not NOT_475(G3117,G2894);
  nand NAND2_39(G3118,G2894,G1503);
  not NOT_476(G3119,G2897);
  nand NAND2_40(G3120,G2897,G1504);
  not NOT_477(G3121,G2900);
  nand NAND2_41(G3122,G2900,G1505);
  not NOT_478(G3123,G2903);
  nand NAND2_42(G3124,G2903,G1506);
  not NOT_479(G3125,G2906);
  nand NAND2_43(G3126,G2906,G1507);
  not NOT_480(G3127,G2909);
  nand NAND2_44(G3128,G2909,G1508);
  not NOT_481(G3129,G2912);
  nand NAND2_45(G3130,G2912,G1509);
  not NOT_482(G3131,G2915);
  nand NAND2_46(G3132,G2918,G1511);
  not NOT_483(G3133,G2918);
  nand NAND2_47(G3134,G2921,G1512);
  not NOT_484(G3135,G2921);
  nand NAND2_48(G3136,G2924,G1513);
  not NOT_485(G3137,G2924);
  nand NAND2_49(G3138,G2927,G1514);
  not NOT_486(G3139,G2927);
  nand NAND2_50(G3140,G2930,G1515);
  not NOT_487(G3141,G2930);
  nand NAND2_51(G3142,G2933,G1516);
  not NOT_488(G3143,G2933);
  nand NAND2_52(G3144,G2936,G1517);
  not NOT_489(G3145,G2936);
  nand NAND2_53(G3146,G2939,G1518);
  not NOT_490(G3147,G2939);
  nand NAND2_54(G3148,G2942,G1519);
  not NOT_491(G3149,G2942);
  not NOT_492(G3150,G2951);
  nand NAND2_55(G3151,G2951,G1582);
  not NOT_493(G3152,G2954);
  nand NAND2_56(G3153,G2954,G1583);
  not NOT_494(G3154,G2957);
  nand NAND2_57(G3155,G2957,G1584);
  nand NAND2_58(G3156,G1377,G3056);
  not NOT_495(G3157,G2960);
  nand NAND2_59(G3158,G2960,G1586);
  not NOT_496(G3159,G2963);
  nand NAND2_60(G3160,G2963,G1587);
  and AND2_202(G3161,G2759,G2774);
  and AND2_203(G3162,G2759,G2774);
  and AND2_204(G3163,G21,G2797);
  not NOT_497(G3164,G2966);
  nand NAND2_61(G3165,G2969,G1589);
  not NOT_498(G3166,G2969);
  nand NAND2_62(G3167,G2972,G1590);
  not NOT_499(G3168,G2972);
  nand NAND2_63(G3169,G1395,G3059);
  nand NAND2_64(G3170,G2975,G1592);
  not NOT_500(G3171,G2975);
  nand NAND2_65(G3172,G2978,G1593);
  not NOT_501(G3173,G2978);
  nand NAND2_66(G3174,G2981,G1594);
  not NOT_502(G3175,G2981);
  and AND2_205(G3176,G2817,G2832);
  and AND2_206(G3177,G2817,G2832);
  not NOT_503(G3178,G2987);
  not NOT_504(G3179,G2990);
  nand NAND2_67(G3180,G2993,G2877);
  not NOT_505(G3181,G2993);
  not NOT_506(G3182,G2996);
  nand NAND2_68(G3183,G2996,G3064);
  not NOT_507(G3184,G3011);
  not NOT_508(G3185,G3014);
  not NOT_509(G3186,G3017);
  not NOT_510(G3187,G3020);
  nand NAND2_69(G3188,G3023,G2878);
  not NOT_511(G3189,G3023);
  nor NOR2_5(G3190,G3065,G2599);
  nor NOR2_6(G3191,G3066,G3067);
  not NOT_512(G3192,G2879);
  nand NAND2_70(G3195,G2629,G3074);
  nand NAND2_71(G3196,G2626,G3075);
  nand NAND2_72(G3197,G2635,G3076);
  nand NAND2_73(G3198,G2632,G3077);
  not NOT_513(G3199,G2883);
  nand NAND2_74(G3202,G2650,G3078);
  nand NAND2_75(G3203,G2647,G3079);
  nand NAND2_76(G3204,G2355,G3080);
  and AND3_191(G3205,G2603,G2332,G3082);
  and AND3_192(G3206,G2328,G2606,G3083);
  and AND3_193(G3207,G3063,G2020,G2031);
  not NOT_514(G3208,G2872);
  not NOT_515(G3211,G2685);
  not NOT_516(G3214,G2945);
  not NOT_517(G3215,G2720);
  not NOT_518(G3218,G2948);
  not NOT_519(G3219,G2744);
  not NOT_520(G3222,G2797);
  not NOT_521(G3225,G2752);
  not NOT_522(G3228,G2752);
  not NOT_523(G3231,G2759);
  not NOT_524(G3234,G2759);
  not NOT_525(G3237,G2780);
  not NOT_526(G3240,G2984);
  not NOT_527(G3241,G2810);
  not NOT_528(G3244,G2817);
  not NOT_529(G3247,G2837);
  not NOT_530(G3250,G2810);
  not NOT_531(G3253,G2817);
  not NOT_532(G3256,G2865);
  not NOT_533(G3259,G2857);
  not NOT_534(G3262,G2865);
  not NOT_535(G3265,G2999);
  not NOT_536(G3266,G3002);
  not NOT_537(G3267,G3005);
  not NOT_538(G3268,G3008);
  not NOT_539(G3269,G3026);
  not NOT_540(G3270,G3029);
  not NOT_541(G3271,G3032);
  not NOT_542(G3272,G3035);
  nand NAND2_77(G3273,G2641,G3097);
  nand NAND2_78(G3274,G2638,G3098);
  nand NAND2_79(G3275,G2659,G3100);
  nand NAND2_80(G3276,G2656,G3101);
  nand NAND2_81(G3277,G3041,G3102);
  nand NAND2_82(G3280,G2363,G3103);
  not NOT_543(G3281,G3060);
  nand NAND2_83(G3282,G1311,G3113);
  nand NAND2_84(G3283,G1314,G3115);
  nand NAND2_85(G3284,G1317,G3117);
  nand NAND2_86(G3285,G1320,G3119);
  nand NAND2_87(G3286,G1323,G3121);
  nand NAND2_88(G3287,G1326,G3123);
  nand NAND2_89(G3288,G1329,G3125);
  nand NAND2_90(G3289,G1332,G3127);
  nand NAND2_91(G3290,G1335,G3129);
  nand NAND2_92(G3291,G1341,G3133);
  nand NAND2_93(G3292,G1344,G3135);
  nand NAND2_94(G3293,G1347,G3137);
  nand NAND2_95(G3294,G1350,G3139);
  nand NAND2_96(G3295,G1353,G3141);
  nand NAND2_97(G3296,G1356,G3143);
  nand NAND2_98(G3297,G1359,G3145);
  nand NAND2_99(G3298,G1362,G3147);
  nand NAND2_100(G3299,G1365,G3149);
  nand NAND2_101(G3300,G1368,G3150);
  nand NAND2_102(G3301,G1371,G3152);
  nand NAND2_103(G3302,G1374,G3154);
  nand NAND2_104(G3303,G3156,G3057);
  nand NAND2_105(G3313,G1380,G3157);
  nand NAND2_106(G3314,G1383,G3159);
  nand NAND2_107(G3315,G1389,G3166);
  nand NAND2_108(G3316,G1392,G3168);
  nand NAND2_109(G3317,G3058,G3169);
  nand NAND2_110(G3331,G1398,G3171);
  nand NAND2_111(G3332,G1401,G3173);
  nand NAND2_112(G3333,G1404,G3175);
  nand NAND2_113(G3334,G2990,G3178);
  nand NAND2_114(G3335,G2987,G3179);
  nand NAND2_115(G3336,G2517,G3181);
  nand NAND2_116(G3337,G2621,G3182);
  nand NAND2_117(G3338,G3014,G3184);
  nand NAND2_118(G3339,G3011,G3185);
  nand NAND2_119(G3340,G3020,G3186);
  nand NAND2_120(G3341,G3017,G3187);
  nand NAND2_121(G3342,G2520,G3189);
  not NOT_544(G3343,G3094);
  nand NAND2_122(G3344,G3195,G3196);
  nand NAND2_123(G3348,G3197,G3198);
  nand NAND2_124(G3351,G3202,G3203);
  nand NAND2_125(G3355,G3204,G3081);
  nor NOR2_7(G3358,G3205,G3084);
  nor NOR2_8(G3359,G3206,G3085);
  or OR2_60(G3360,G2804,G3163);
  nand NAND2_126(G3363,G3002,G3265);
  nand NAND2_127(G3364,G2999,G3266);
  nand NAND2_128(G3365,G3008,G3267);
  nand NAND2_129(G3366,G3005,G3268);
  nand NAND2_130(G3367,G3029,G3269);
  nand NAND2_131(G3368,G3026,G3270);
  nand NAND2_132(G3369,G3035,G3271);
  nand NAND2_133(G3370,G3032,G3272);
  nand NAND2_134(G3371,G3191,G3190);
  not NOT_545(G3374,G3060);
  nand NAND2_135(G3377,G3273,G3274);
  nand NAND2_136(G3380,G3275,G3276);
  nand NAND2_137(G3383,G3280,G3104);
  nand NAND2_138(G3386,G3282,G3114);
  nand NAND2_139(G3393,G3283,G3116);
  nand NAND2_140(G3404,G3284,G3118);
  nand NAND2_141(G3415,G3285,G3120);
  nand NAND2_142(G3421,G3286,G3122);
  nand NAND2_143(G3428,G3287,G3124);
  nand NAND2_144(G3438,G3288,G3126);
  nand NAND2_145(G3449,G3289,G3128);
  nand NAND2_146(G3459,G3290,G3130);
  not NOT_546(G3466,G3211);
  nand NAND2_147(G3467,G3132,G3291);
  nand NAND2_148(G3474,G3134,G3292);
  nand NAND2_149(G3485,G3136,G3293);
  nand NAND2_150(G3495,G3138,G3294);
  nand NAND2_151(G3503,G3140,G3295);
  nand NAND2_152(G3517,G3142,G3296);
  nand NAND2_153(G3533,G3144,G3297);
  nand NAND2_154(G3546,G3146,G3298);
  nand NAND2_155(G3552,G3148,G3299);
  nand NAND2_156(G3559,G3300,G3151);
  nand NAND2_157(G3570,G3301,G3153);
  nand NAND2_158(G3576,G3302,G3155);
  nand NAND2_159(G3583,G3313,G3158);
  nand NAND2_160(G3594,G3314,G3160);
  nand NAND2_161(G3604,G3222,G1588);
  not NOT_547(G3605,G3222);
  not NOT_548(G3606,G3225);
  not NOT_549(G3607,G3228);
  not NOT_550(G3608,G3231);
  not NOT_551(G3609,G3234);
  not NOT_552(G3610,G3237);
  nand NAND2_162(G3611,G3165,G3315);
  nand NAND2_163(G3621,G3167,G3316);
  nand NAND2_164(G3629,G3170,G3331);
  nand NAND2_165(G3645,G3172,G3332);
  nand NAND2_166(G3658,G3174,G3333);
  not NOT_553(G3664,G3244);
  not NOT_554(G3665,G3253);
  nand NAND2_167(G3666,G3334,G3335);
  nand NAND2_168(G3670,G3180,G3336);
  nand NAND2_169(G3674,G3337,G3183);
  nand NAND2_170(G3677,G3338,G3339);
  nand NAND2_171(G3681,G3340,G3341);
  nand NAND2_172(G3685,G3188,G3342);
  and AND2_207(G3688,G3208,G2872);
  not NOT_555(G3689,G3215);
  not NOT_556(G3690,G3219);
  not NOT_557(G3691,G3241);
  not NOT_558(G3692,G3247);
  not NOT_559(G3693,G3250);
  not NOT_560(G3694,G3256);
  not NOT_561(G3695,G3259);
  not NOT_562(G3696,G3262);
  nand NAND2_173(G3697,G3365,G3366);
  nand NAND2_174(G3700,G3363,G3364);
  nand NAND2_175(G3703,G3369,G3370);
  nand NAND2_176(G3706,G3367,G3368);
  not NOT_563(G3709,G3277);
  nand NAND2_177(G3710,G3359,G3358);
  and AND2_208(G3713,G3303,G2788);
  nand NAND2_178(G3714,G1386,G3605);
  not NOT_564(G3715,G3360);
  and AND2_209(G3716,G3317,G2844);
  and AND2_210(G3717,G3317,G2844);
  not NOT_565(G3718,G3371);
  nand NAND2_179(G3719,G3371,G3343);
  not NOT_566(G3720,G3344);
  not NOT_567(G3723,G3351);
  not NOT_568(G3726,G3348);
  not NOT_569(G3729,G3348);
  not NOT_570(G3732,G3355);
  not NOT_571(G3735,G3355);
  not NOT_572(G3738,G3383);
  or OR2_61(G3739,G3208,G3688);
  not NOT_573(G3742,G3303);
  not NOT_574(G3745,G3317);
  not NOT_575(G3748,G3317);
  not NOT_576(G3751,G3374);
  nand NAND2_180(G3752,G3374,G3099);
  not NOT_577(G3753,G3377);
  not NOT_578(G3754,G3380);
  nand NAND2_181(G3755,G3380,G3709);
  and AND2_211(G3756,G3467,G2711);
  and AND3_194(G3757,G3474,G3467,G2715);
  and AND4_5(G3758,G3485,G3467,G2720,G3474);
  and AND4_6(G3759,G3559,G2752,G2780,G2759);
  and AND2_212(G3760,G3386,G2675);
  and AND3_195(G3761,G3393,G3386,G2679);
  and AND4_7(G3762,G3404,G3386,G2685,G3393);
  and AND4_8(G3763,G3611,G2810,G2837,G2817);
  not NOT_579(G3764,G3415);
  and AND4_9(G3765,G3393,G3415,G3404,G3386);
  and AND2_213(G3768,G3393,G2679);
  and AND3_196(G3769,G3404,G2685,G3393);
  and AND3_197(G3770,G3415,G3404,G3393);
  and AND2_214(G3771,G3393,G2679);
  and AND3_198(G3772,G2685,G3404,G3393);
  and AND2_215(G3773,G3404,G2685);
  and AND2_216(G3774,G3415,G3404);
  and AND2_217(G3775,G3404,G2685);
  and AND5_0(G3776,G3428,G3459,G3438,G3421,G3449);
  and AND2_218(G3779,G3421,G2693);
  and AND3_199(G3780,G3428,G3421,G2696);
  and AND4_10(G3781,G3438,G3421,G2700,G3428);
  and AND5_1(G3782,G3449,G3438,G3421,G2705,G3428);
  and AND2_219(G3783,G3428,G2696);
  and AND3_200(G3784,G3438,G2700,G3428);
  and AND4_11(G3785,G3449,G3438,G2705,G3428);
  and AND5_2(G3786,G2,G3459,G3438,G3449,G3428);
  and AND2_220(G3787,G2700,G3438);
  and AND3_201(G3788,G3449,G3438,G2705);
  and AND4_12(G3789,G2,G3459,G3438,G3449);
  and AND2_221(G3790,G3449,G2705);
  and AND3_202(G3791,G2,G3459,G3449);
  and AND2_222(G3792,G2,G3459);
  and AND4_13(G3793,G3546,G3485,G3474,G3467);
  and AND2_223(G3796,G3474,G2715);
  and AND3_203(G3797,G3485,G2720,G3474);
  and AND3_204(G3798,G3546,G3485,G3474);
  and AND2_224(G3799,G3474,G2715);
  and AND3_205(G3800,G3485,G2720,G3474);
  and AND2_225(G3801,G3485,G2720);
  and AND5_3(G3802,G3552,G3533,G3517,G3503,G3495);
  and AND2_226(G3805,G3495,G2727);
  and AND3_206(G3806,G3503,G3495,G2731);
  and AND4_14(G3807,G3517,G3495,G2737,G3503);
  and AND5_4(G3808,G3533,G3517,G3495,G2744,G3503);
  and AND2_227(G3809,G3503,G2731);
  and AND3_207(G3810,G3517,G2737,G3503);
  and AND4_15(G3811,G3533,G3517,G2744,G3503);
  and AND4_16(G3812,G3552,G3517,G3503,G3533);
  and AND2_228(G3813,G3503,G2731);
  and AND3_208(G3814,G3517,G2737,G3503);
  and AND4_17(G3815,G3533,G3517,G2744,G3503);
  and AND2_229(G3816,G3517,G2737);
  and AND3_209(G3817,G3533,G3517,G2744);
  and AND3_210(G3818,G3552,G3517,G3533);
  and AND2_230(G3819,G3517,G2737);
  and AND3_211(G3820,G3533,G3517,G2744);
  and AND2_231(G3821,G3533,G2744);
  and AND2_232(G3822,G3546,G3485);
  and AND2_233(G3823,G3552,G3533);
  not NOT_580(G3824,G3570);
  and AND4_18(G3825,G2759,G3570,G3559,G2752);
  and AND3_212(G3828,G3559,G2780,G2759);
  and AND3_213(G3829,G3570,G3559,G2759);
  and AND3_214(G3830,G2780,G3559,G2759);
  and AND2_234(G3831,G3559,G2780);
  and AND2_235(G3832,G3570,G3559);
  and AND2_236(G3833,G3559,G2780);
  and AND5_5(G3834,G3303,G2797,G3583,G3576,G3594);
  and AND2_237(G3837,G3576,G2540);
  and AND3_215(G3838,G3303,G3576,G2788);
  and AND4_19(G3839,G3583,G3576,G2792,G3303);
  and AND5_6(G3840,G3594,G3583,G3576,G2804,G3303);
  and AND3_216(G3841,G3583,G2792,G3303);
  and AND4_20(G3842,G3594,G3583,G2804,G3303);
  and AND5_7(G3843,G21,G2797,G3583,G3594,G3303);
  and AND2_238(G3844,G2792,G3583);
  and AND3_217(G3845,G3594,G3583,G2804);
  and AND4_21(G3846,G21,G2797,G3583,G3594);
  and AND2_239(G3847,G3594,G2804);
  and AND3_218(G3848,G21,G2797,G3594);
  nand NAND2_182(G3849,G3604,G3714);
  and AND4_22(G3852,G3658,G3611,G2817,G2810);
  and AND3_219(G3855,G3611,G2837,G2817);
  and AND3_220(G3856,G3658,G3611,G2817);
  and AND3_221(G3857,G3611,G2837,G2817);
  and AND2_240(G3858,G3611,G2837);
  and AND5_8(G3859,G2865,G3645,G3629,G3317,G3621);
  and AND2_241(G3862,G3621,G2543);
  and AND3_222(G3863,G3317,G3621,G2844);
  and AND4_23(G3864,G3629,G3621,G2850,G3317);
  and AND5_9(G3865,G3645,G3629,G3621,G2857,G3317);
  and AND3_223(G3866,G3629,G2850,G3317);
  and AND4_24(G3867,G3645,G3629,G2857,G3317);
  and AND4_25(G3868,G2865,G3629,G3317,G3645);
  and AND3_224(G3869,G3629,G2850,G3317);
  and AND4_26(G3870,G3645,G3629,G2857,G3317);
  and AND2_242(G3871,G3629,G2850);
  and AND3_225(G3872,G3645,G3629,G2857);
  and AND3_226(G3873,G2865,G3629,G3645);
  and AND2_243(G3874,G3629,G2850);
  and AND3_227(G3875,G3645,G3629,G2857);
  and AND2_244(G3876,G3645,G2857);
  and AND2_245(G3877,G3658,G3611);
  and AND2_246(G3878,G2865,G3645);
  not NOT_581(G3879,G3666);
  not NOT_582(G3882,G3670);
  not NOT_583(G3885,G3677);
  not NOT_584(G3888,G3681);
  not NOT_585(G3891,G3674);
  not NOT_586(G3894,G3674);
  not NOT_587(G3897,G3685);
  not NOT_588(G3900,G3685);
  nand NAND2_183(G3903,G3094,G3718);
  not NOT_589(G3904,G3710);
  nand NAND2_184(G3905,G3710,G3738);
  not NOT_590(G3906,G3459);
  not NOT_591(G3909,G3386);
  not NOT_592(G3912,G3386);
  not NOT_593(G3915,G3393);
  not NOT_594(G3918,G3393);
  not NOT_595(G3921,G3404);
  not NOT_596(G3924,G3404);
  not NOT_597(G3927,G3421);
  not NOT_598(G3930,G3428);
  not NOT_599(G3933,G3438);
  not NOT_600(G3936,G3449);
  not NOT_601(G3939,G3546);
  not NOT_602(G3942,G3485);
  not NOT_603(G3945,G3467);
  not NOT_604(G3948,G3474);
  not NOT_605(G3951,G3546);
  not NOT_606(G3954,G3485);
  not NOT_607(G3957,G3467);
  not NOT_608(G3960,G3474);
  not NOT_609(G3963,G3552);
  not NOT_610(G3966,G3533);
  not NOT_611(G3969,G3495);
  not NOT_612(G3972,G3517);
  not NOT_613(G3975,G3503);
  not NOT_614(G3978,G3503);
  not NOT_615(G3981,G3552);
  not NOT_616(G3984,G3533);
  not NOT_617(G3987,G3495);
  not NOT_618(G3990,G3517);
  not NOT_619(G3993,G3559);
  not NOT_620(G3996,G3559);
  not NOT_621(G3999,G3576);
  not NOT_622(G4002,G3583);
  not NOT_623(G4005,G3594);
  not NOT_624(G4008,G3658);
  not NOT_625(G4011,G3611);
  not NOT_626(G4014,G3658);
  not NOT_627(G4017,G3611);
  not NOT_628(G4020,G3645);
  not NOT_629(G4023,G3621);
  not NOT_630(G4026,G3629);
  not NOT_631(G4029,G3645);
  not NOT_632(G4032,G3621);
  not NOT_633(G4035,G3629);
  not NOT_634(G4038,G3697);
  not NOT_635(G4039,G3700);
  not NOT_636(G4040,G3703);
  not NOT_637(G4041,G3706);
  nand NAND2_185(G4042,G2644,G3751);
  nand NAND2_186(G4043,G3277,G3754);
  or OR4_4(G4044,G2667,G3756,G3757,G3758);
  or OR4_5(G4045,G2492,G3109,G3110,G3759);
  or OR4_6(G4046,G2670,G3760,G3761,G3762);
  or OR4_7(G4047,G2492,G3111,G3112,G3763);
  or OR5_0(G4048,G2692,G3779,G3780,G3781,G3782);
  or OR2_62(G4051,G2715,G3801);
  or OR5_1(G4054,G2726,G3805,G3806,G3807,G3808);
  or OR2_63(G4058,G2737,G3821);
  or OR5_2(G4061,G2787,G3837,G3838,G3839,G3840);
  not NOT_638(G4064,G3742);
  or OR2_64(G4065,G2832,G3858);
  or OR5_3(G4068,G2843,G3862,G3863,G3864,G3865);
  or OR2_65(G4072,G2850,G3876);
  not NOT_639(G4075,G3745);
  not NOT_640(G4076,G3748);
  nand NAND2_187(G4077,G3903,G3719);
  not NOT_641(G4080,G3726);
  not NOT_642(G4081,G3729);
  not NOT_643(G4082,G3732);
  not NOT_644(G4083,G3735);
  and AND3_228(G4084,G3344,G2879,G3726);
  and AND3_229(G4085,G3720,G3192,G3729);
  and AND3_230(G4086,G3351,G2883,G3732);
  and AND3_231(G4087,G3723,G3199,G3735);
  nand NAND2_188(G4088,G3383,G3904);
  nand NAND2_189(G4089,G3739,G61);
  or OR4_8(G4092,G2675,G3768,G3769,G3770);
  nor NOR3_0(G4095,G2675,G3771,G3772);
  or OR3_28(G4098,G2679,G3773,G3774);
  nor NOR2_9(G4101,G2679,G3775);
  or OR5_4(G4104,G2693,G3783,G3784,G3785,G3786);
  or OR4_9(G4107,G2696,G3787,G3788,G3789);
  or OR3_29(G4110,G2700,G3790,G3791);
  or OR2_66(G4113,G2705,G3792);
  or OR4_10(G4116,G2711,G3796,G3797,G3798);
  nor NOR3_1(G4119,G2711,G3799,G3800);
  or OR4_11(G4122,G2731,G3816,G3817,G3818);
  or OR5_5(G4125,G2727,G3809,G3810,G3811,G3812);
  nor NOR3_2(G4128,G2731,G3819,G3820);
  nor NOR4_0(G4131,G2727,G3813,G3814,G3815);
  or OR4_12(G4134,G2770,G3161,G3828,G3829);
  nor NOR3_3(G4137,G2770,G3162,G3830);
  or OR3_30(G4140,G2774,G3831,G3832);
  nor NOR2_10(G4143,G2774,G3833);
  or OR5_6(G4146,G2540,G3713,G3841,G3842,G3843);
  or OR4_13(G4149,G2788,G3844,G3845,G3846);
  or OR3_31(G4152,G2792,G3847,G3848);
  or OR4_14(G4155,G2828,G3176,G3855,G3856);
  nor NOR3_4(G4158,G2828,G3177,G3857);
  or OR4_15(G4161,G2844,G3871,G3872,G3873);
  or OR5_7(G4164,G2543,G3716,G3866,G3867,G3868);
  nor NOR3_5(G4167,G2844,G3874,G3875);
  nor NOR4_1(G4170,G2543,G3717,G3869,G3870);
  nand NAND2_190(G4173,G3700,G4038);
  nand NAND2_191(G4174,G3697,G4039);
  nand NAND2_192(G4175,G3706,G4040);
  nand NAND2_193(G4176,G3703,G4041);
  nand NAND2_194(G4177,G4042,G3752);
  nand NAND2_195(G4180,G3755,G4043);
  not NOT_645(G4183,G3849);
  nand NAND2_196(G4184,G3906,G1510);
  not NOT_646(G4185,G3906);
  not NOT_647(G4186,G3909);
  not NOT_648(G4187,G3912);
  not NOT_649(G4188,G3915);
  not NOT_650(G4189,G3918);
  nand NAND2_197(G4190,G3921,G3131);
  not NOT_651(G4191,G3921);
  nand NAND2_198(G4192,G3924,G3466);
  not NOT_652(G4193,G3924);
  and AND2_247(G4194,G3776,G2);
  not NOT_653(G4195,G3927);
  not NOT_654(G4196,G3930);
  not NOT_655(G4197,G3933);
  not NOT_656(G4198,G3936);
  not NOT_657(G4199,G3802);
  not NOT_658(G4200,G3948);
  not NOT_659(G4201,G3960);
  not NOT_660(G4202,G3975);
  not NOT_661(G4203,G3978);
  nand NAND2_199(G4204,G3993,G3164);
  not NOT_662(G4205,G3993);
  nand NAND2_200(G4206,G3996,G3610);
  not NOT_663(G4207,G3996);
  and AND2_248(G4208,G3834,G21);
  not NOT_664(G4209,G3999);
  not NOT_665(G4210,G4002);
  nand NAND2_201(G4211,G4005,G3715);
  not NOT_666(G4212,G4005);
  not NOT_667(G4213,G3859);
  not NOT_668(G4214,G3891);
  not NOT_669(G4215,G3894);
  not NOT_670(G4216,G3897);
  not NOT_671(G4217,G3900);
  and AND3_232(G4218,G3670,G3666,G3891);
  and AND3_233(G4219,G3882,G3879,G3894);
  and AND3_234(G4220,G3681,G3677,G3897);
  and AND3_235(G4221,G3888,G3885,G3900);
  and AND3_236(G4222,G3849,G1264,G2003);
  and AND3_237(G4223,G3192,G3344,G4080);
  and AND3_238(G4224,G2879,G3720,G4081);
  and AND3_239(G4225,G3199,G3351,G4082);
  and AND3_240(G4226,G2883,G3723,G4083);
  nand NAND2_202(G4227,G4088,G3905);
  not NOT_672(G4230,G3939);
  not NOT_673(G4231,G3942);
  not NOT_674(G4232,G3945);
  not NOT_675(G4233,G3951);
  not NOT_676(G4234,G3954);
  not NOT_677(G4235,G3957);
  not NOT_678(G4236,G3963);
  not NOT_679(G4237,G3966);
  not NOT_680(G4238,G3969);
  not NOT_681(G4239,G3972);
  not NOT_682(G4240,G3990);
  not NOT_683(G4241,G3981);
  not NOT_684(G4242,G3984);
  not NOT_685(G4243,G3987);
  not NOT_686(G4244,G4008);
  not NOT_687(G4245,G4011);
  not NOT_688(G4246,G4014);
  not NOT_689(G4247,G4017);
  not NOT_690(G4248,G4020);
  not NOT_691(G4249,G4023);
  not NOT_692(G4250,G4026);
  not NOT_693(G4251,G4035);
  not NOT_694(G4252,G4029);
  not NOT_695(G4253,G4032);
  nand NAND2_203(G4254,G4173,G4174);
  nand NAND2_204(G4257,G4175,G4176);
  and AND2_249(G4260,G3793,G4054);
  and AND2_250(G4261,G4061,G3825);
  and AND2_251(G4262,G4048,G3765);
  and AND2_252(G4263,G3852,G4068);
  not NOT_696(G4264,G4077);
  nand NAND2_205(G4265,G1338,G4185);
  not NOT_697(G4266,G4092);
  nand NAND2_206(G4267,G4092,G4186);
  not NOT_698(G4268,G4095);
  nand NAND2_207(G4269,G4095,G4187);
  not NOT_699(G4270,G4098);
  nand NAND2_208(G4271,G4098,G4188);
  not NOT_700(G4272,G4101);
  nand NAND2_209(G4273,G4101,G4189);
  nand NAND2_210(G4274,G2915,G4191);
  nand NAND2_211(G4275,G3211,G4193);
  or OR2_67(G4276,G4048,G4194);
  not NOT_701(G4282,G4104);
  nand NAND2_212(G4283,G4104,G4195);
  not NOT_702(G4284,G4107);
  nand NAND2_213(G4285,G4107,G4196);
  not NOT_703(G4286,G4110);
  nand NAND2_214(G4287,G4110,G4197);
  not NOT_704(G4288,G4113);
  nand NAND2_215(G4289,G4113,G4198);
  not NOT_705(G4290,G4054);
  not NOT_706(G4293,G4134);
  nand NAND2_216(G4294,G4134,G3606);
  not NOT_707(G4295,G4137);
  nand NAND2_217(G4296,G4137,G3607);
  not NOT_708(G4297,G4140);
  nand NAND2_218(G4298,G4140,G3608);
  not NOT_709(G4299,G4143);
  nand NAND2_219(G4300,G4143,G3609);
  nand NAND2_220(G4301,G2966,G4205);
  nand NAND2_221(G4302,G3237,G4207);
  or OR2_68(G4303,G4061,G4208);
  not NOT_710(G4309,G4146);
  nand NAND2_222(G4310,G4146,G4209);
  not NOT_711(G4311,G4149);
  nand NAND2_223(G4312,G4149,G4064);
  not NOT_712(G4313,G4152);
  nand NAND2_224(G4314,G4152,G4210);
  nand NAND2_225(G4315,G3360,G4212);
  not NOT_713(G4316,G4068);
  and AND3_241(G4319,G3879,G3670,G4214);
  and AND3_242(G4320,G3666,G3882,G4215);
  and AND3_243(G4321,G3885,G3681,G4216);
  and AND3_244(G4322,G3677,G3888,G4217);
  or OR3_32(G4323,G2600,G4222,G2324);
  nor NOR2_11(G4329,G4223,G4084);
  nor NOR2_12(G4330,G4224,G4085);
  nor NOR2_13(G4331,G4225,G4086);
  nor NOR2_14(G4332,G4226,G4087);
  not NOT_714(G4333,G4180);
  and AND2_253(G4334,G3739,G4089);
  and AND2_254(G4335,G4089,G61);
  or OR2_69(G4336,G4051,G3822);
  not NOT_715(G4339,G4116);
  not NOT_716(G4340,G4051);
  not NOT_717(G4343,G4119);
  not NOT_718(G4344,G4122);
  nand NAND2_226(G4345,G4122,G3218);
  or OR2_70(G4346,G4058,G3823);
  not NOT_719(G4349,G4125);
  not NOT_720(G4350,G4128);
  nand NAND2_227(G4351,G4128,G3690);
  not NOT_721(G4352,G4058);
  not NOT_722(G4355,G4131);
  or OR2_71(G4356,G4065,G3877);
  not NOT_723(G4359,G4155);
  not NOT_724(G4360,G4065);
  not NOT_725(G4363,G4158);
  or OR2_72(G4364,G4072,G3878);
  not NOT_726(G4367,G4161);
  not NOT_727(G4368,G4164);
  not NOT_728(G4369,G4167);
  nand NAND2_228(G4370,G4167,G3695);
  not NOT_729(G4371,G4072);
  not NOT_730(G4374,G4170);
  not NOT_731(G4375,G4177);
  nand NAND2_229(G4376,G4177,G3753);
  not NOT_732(G4377,G4227);
  nand NAND2_230(G4378,G4184,G4265);
  nand NAND2_231(G4381,G3909,G4266);
  nand NAND2_232(G4382,G3912,G4268);
  nand NAND2_233(G4383,G3915,G4270);
  nand NAND2_234(G4384,G3918,G4272);
  nand NAND2_235(G4385,G4190,G4274);
  nand NAND2_236(G4386,G4192,G4275);
  nand NAND2_237(G4387,G3927,G4282);
  nand NAND2_238(G4388,G3930,G4284);
  nand NAND2_239(G4389,G3933,G4286);
  nand NAND2_240(G4390,G3936,G4288);
  nand NAND2_241(G4391,G3225,G4293);
  nand NAND2_242(G4392,G3228,G4295);
  nand NAND2_243(G4393,G3231,G4297);
  nand NAND2_244(G4394,G3234,G4299);
  nand NAND2_245(G4395,G4204,G4301);
  nand NAND2_246(G4396,G4206,G4302);
  nand NAND2_247(G4397,G3999,G4309);
  nand NAND2_248(G4398,G3742,G4311);
  nand NAND2_249(G4399,G4002,G4313);
  nand NAND2_250(G4400,G4211,G4315);
  nor NOR2_15(G4403,G4319,G4218);
  nor NOR2_16(G4404,G4320,G4219);
  nor NOR2_17(G4405,G4321,G4220);
  nor NOR2_18(G4406,G4322,G4221);
  not NOT_733(G4407,G4254);
  not NOT_734(G4408,G4257);
  or OR2_73(G4409,G4334,G4335);
  nand NAND2_251(G4413,G2948,G4344);
  nand NAND2_252(G4414,G3219,G4350);
  nand NAND2_253(G4415,G3259,G4369);
  nand NAND2_254(G4416,G3377,G4375);
  nand NAND2_255(G4417,G4330,G4329);
  nand NAND2_256(G4420,G4332,G4331);
  and AND3_245(G4423,G4323,G1554,G1565);
  and AND3_246(G4424,G4323,G1629,G1640);
  and AND3_247(G4425,G4323,G1652,G1663);
  and AND3_248(G4426,G4323,G1674,G1685);
  nand NAND2_257(G4427,G4381,G4267);
  nand NAND2_258(G4428,G4382,G4269);
  nand NAND2_259(G4429,G4383,G4271);
  nand NAND2_260(G4430,G4384,G4273);
  not NOT_735(G4431,G4385);
  not NOT_736(G4432,G4276);
  nand NAND2_261(G4437,G4387,G4283);
  nand NAND2_262(G4440,G4388,G4285);
  nand NAND2_263(G4443,G4389,G4287);
  nand NAND2_264(G4446,G4390,G4289);
  and AND2_255(G4449,G4276,G3764);
  and AND2_256(G4450,G4290,G4199);
  nand NAND2_265(G4453,G4391,G4294);
  nand NAND2_266(G4454,G4392,G4296);
  nand NAND2_267(G4455,G4393,G4298);
  nand NAND2_268(G4456,G4394,G4300);
  not NOT_737(G4457,G4395);
  not NOT_738(G4458,G4303);
  nand NAND2_269(G4463,G4397,G4310);
  nand NAND2_270(G4466,G4398,G4312);
  nand NAND2_271(G4469,G4399,G4314);
  and AND2_257(G4472,G4303,G3824);
  and AND2_258(G4473,G4316,G4213);
  not NOT_739(G4476,G4336);
  nand NAND2_272(G4477,G4336,G3214);
  not NOT_740(G4478,G4340);
  nand NAND2_273(G4479,G4340,G3689);
  nand NAND2_274(G4480,G4345,G4413);
  not NOT_741(G4483,G4346);
  nand NAND2_275(G4484,G4351,G4414);
  not NOT_742(G4487,G4352);
  not NOT_743(G4488,G4356);
  nand NAND2_276(G4489,G4356,G3240);
  not NOT_744(G4490,G4360);
  nand NAND2_277(G4491,G4360,G3692);
  not NOT_745(G4492,G4364);
  nand NAND2_278(G4493,G4364,G4367);
  nand NAND2_279(G4494,G4370,G4415);
  not NOT_746(G4497,G4371);
  nand NAND2_280(G4498,G4404,G4403);
  nand NAND2_281(G4501,G4406,G4405);
  nand NAND2_282(G4504,G4416,G4376);
  not NOT_747(G4507,G4378);
  not NOT_748(G4508,G4400);
  and AND3_249(G4509,G4409,G171,G1242);
  not NOT_749(G4510,G4428);
  not NOT_750(G4511,G4430);
  and AND2_259(G4512,G4276,G4427);
  and AND2_260(G4513,G4276,G4429);
  and AND2_261(G4514,G4276,G4431);
  not NOT_751(G4515,G4454);
  not NOT_752(G4516,G4456);
  and AND2_262(G4517,G4303,G4453);
  and AND2_263(G4518,G4303,G4455);
  and AND2_264(G4519,G4303,G4457);
  and AND3_250(G4520,G4378,G1248,G1981);
  and AND3_251(G4521,G4400,G1264,G2003);
  not NOT_753(G4522,G4417);
  not NOT_754(G4523,G4420);
  nand NAND2_283(G4524,G4420,G4333);
  nand NAND2_284(G4525,G2945,G4476);
  nand NAND2_285(G4526,G3215,G4478);
  nand NAND2_286(G4527,G2984,G4488);
  nand NAND2_287(G4528,G3247,G4490);
  nand NAND2_288(G4529,G4161,G4492);
  not NOT_755(G4530,G4446);
  not NOT_756(G4531,G4443);
  not NOT_757(G4532,G4440);
  not NOT_758(G4533,G4437);
  not NOT_759(G4534,G4469);
  not NOT_760(G4535,G4466);
  not NOT_761(G4536,G4463);
  and AND2_265(G4537,G4510,G4432);
  and AND2_266(G4538,G4511,G4432);
  and AND2_267(G4539,G4386,G4432);
  and AND2_268(G4540,G3415,G4432);
  not NOT_762(G4541,G4450);
  and AND2_269(G4542,G4515,G4458);
  and AND2_270(G4543,G4516,G4458);
  and AND2_271(G4544,G4396,G4458);
  and AND2_272(G4545,G3570,G4458);
  not NOT_763(G4546,G4473);
  not NOT_764(G4547,G4498);
  nand NAND2_289(G4548,G4498,G4407);
  not NOT_765(G4549,G4501);
  nand NAND2_290(G4550,G4501,G4408);
  and AND3_252(G4551,G4446,G1248,G1981);
  and AND3_253(G4552,G4443,G1248,G1981);
  and AND3_254(G4553,G4440,G1248,G1981);
  or OR3_33(G4554,G3068,G4520,G2320);
  and AND3_255(G4560,G4469,G1264,G2003);
  and AND3_256(G4561,G4466,G1264,G2003);
  or OR3_34(G4562,G3072,G4521,G2325);
  nand NAND2_291(G4568,G4504,G4522);
  not NOT_766(G4569,G4504);
  nand NAND2_292(G4570,G4180,G4523);
  and AND3_257(G4571,G4437,G1280,G2031);
  and AND3_258(G4572,G4463,G1294,G2053);
  nand NAND2_293(G4573,G4477,G4525);
  nand NAND2_294(G4576,G4479,G4526);
  not NOT_767(G4579,G4480);
  nand NAND2_295(G4580,G4480,G4483);
  not NOT_768(G4581,G4484);
  nand NAND2_296(G4582,G4484,G4487);
  nand NAND2_297(G4583,G4489,G4527);
  nand NAND2_298(G4586,G4491,G4528);
  nand NAND2_299(G4589,G4493,G4529);
  not NOT_769(G4592,G4494);
  nand NAND2_300(G4593,G4494,G4497);
  or OR2_74(G4594,G4537,G4512);
  or OR2_75(G4597,G4538,G4513);
  or OR2_76(G4600,G4539,G4514);
  or OR2_77(G4603,G4540,G4449);
  or OR2_78(G4606,G4542,G4517);
  or OR2_79(G4613,G4543,G4518);
  or OR2_80(G4616,G4544,G4519);
  or OR2_81(G4619,G4545,G4472);
  nand NAND2_301(G4622,G4254,G4547);
  nand NAND2_302(G4623,G4257,G4549);
  or OR3_35(G4624,G3069,G4551,G2321);
  or OR3_36(G4630,G3070,G4552,G2322);
  or OR3_37(G4636,G3071,G4553,G2323);
  or OR3_38(G4642,G3073,G4560,G2326);
  or OR3_39(G4648,G2516,G4561,G2327);
  nand NAND2_303(G4654,G4417,G4569);
  nand NAND2_304(G4655,G4570,G4524);
  or OR3_40(G4658,G3086,G4571,G2339);
  or OR3_41(G4664,G3090,G4572,G2344);
  nand NAND2_305(G4670,G4346,G4579);
  nand NAND2_306(G4671,G4352,G4581);
  nand NAND2_307(G4672,G4371,G4592);
  and AND3_259(G4673,G4554,G718,G1565);
  and AND3_260(G4674,G4562,G1554,G1565);
  and AND3_261(G4675,G4554,G780,G1640);
  and AND3_262(G4676,G4562,G1629,G1640);
  and AND3_263(G4677,G4554,G860,G1663);
  and AND3_264(G4678,G4562,G1652,G1663);
  and AND3_265(G4679,G4562,G1674,G1685);
  and AND3_266(G4680,G4554,G884,G1685);
  nand NAND2_308(G4681,G4622,G4548);
  nand NAND2_309(G4684,G4623,G4550);
  nand NAND2_310(G4687,G4568,G4654);
  not NOT_770(G4690,G4573);
  nand NAND2_311(G4691,G4573,G4339);
  not NOT_771(G4692,G4576);
  nand NAND2_312(G4693,G4576,G4343);
  nand NAND2_313(G4694,G4670,G4580);
  nand NAND2_314(G4697,G4671,G4582);
  not NOT_772(G4700,G4583);
  nand NAND2_315(G4701,G4583,G4359);
  not NOT_773(G4702,G4586);
  nand NAND2_316(G4703,G4586,G4363);
  not NOT_774(G4704,G4589);
  nand NAND2_317(G4705,G4589,G4368);
  nand NAND2_318(G4706,G4672,G4593);
  not NOT_775(G4709,G4603);
  not NOT_776(G4710,G4600);
  not NOT_777(G4711,G4597);
  not NOT_778(G4712,G4594);
  not NOT_779(G4713,G4619);
  not NOT_780(G4714,G4616);
  not NOT_781(G4715,G4613);
  not NOT_782(G4716,G4606);
  and AND3_267(G4717,G4664,G1526,G1537);
  and AND3_268(G4718,G4658,G694,G1537);
  or OR4_16(G4719,G4423,G4673,G2162,G1465);
  and AND3_269(G4720,G4624,G718,G1565);
  and AND3_270(G4721,G4642,G1554,G1565);
  and AND3_271(G4722,G4630,G718,G1565);
  and AND3_272(G4723,G4648,G1554,G1565);
  and AND3_273(G4724,G4636,G718,G1565);
  and AND3_274(G4725,G4664,G1601,G1612);
  and AND3_275(G4726,G4658,G756,G1612);
  or OR4_17(G4727,G4424,G4675,G2173,G1474);
  and AND3_276(G4728,G4624,G780,G1640);
  and AND3_277(G4729,G4642,G1629,G1640);
  and AND3_278(G4730,G4630,G780,G1640);
  and AND3_279(G4731,G4648,G1629,G1640);
  and AND3_280(G4732,G4636,G780,G1640);
  and AND3_281(G4733,G4664,G1914,G1925);
  and AND3_282(G4734,G4658,G1184,G1925);
  and AND3_283(G4735,G4648,G1652,G1663);
  and AND3_284(G4736,G4636,G860,G1663);
  and AND3_285(G4737,G4642,G1652,G1663);
  and AND3_286(G4738,G4630,G860,G1663);
  and AND3_287(G4739,G4624,G860,G1663);
  and AND3_288(G4740,G4664,G1948,G1959);
  and AND3_289(G4741,G4658,G1218,G1959);
  and AND3_290(G4742,G4648,G1674,G1685);
  and AND3_291(G4743,G4636,G884,G1685);
  and AND3_292(G4744,G4642,G1674,G1685);
  and AND3_293(G4745,G4630,G884,G1685);
  and AND3_294(G4746,G4624,G884,G1685);
  and AND3_295(G4747,G4606,G171,G170);
  not NOT_783(G4748,G4655);
  and AND2_273(G4749,G4655,G1941);
  and AND3_296(G4750,G4603,G1280,G2031);
  and AND3_297(G4751,G4600,G1280,G2031);
  and AND3_298(G4752,G4597,G1280,G2031);
  and AND3_299(G4753,G4594,G1280,G2031);
  and AND3_300(G4754,G4619,G1294,G2053);
  and AND3_301(G4755,G4616,G1294,G2053);
  and AND3_302(G4756,G4613,G1294,G2053);
  and AND3_303(G4757,G4606,G1294,G2053);
  nand NAND2_319(G4758,G4409,G4606);
  nand NAND2_320(G4761,G4116,G4690);
  nand NAND2_321(G4762,G4119,G4692);
  nand NAND2_322(G4763,G4155,G4700);
  nand NAND2_323(G4764,G4158,G4702);
  nand NAND2_324(G4765,G4164,G4704);
  or OR4_18(G4766,G4717,G4718,G2157,G1460);
  or OR4_19(G4767,G4674,G4720,G2163,G1466);
  or OR4_20(G4768,G4721,G4722,G2164,G1467);
  or OR4_21(G4769,G4723,G4724,G2165,G1468);
  or OR4_22(G4770,G4725,G4726,G2168,G1469);
  or OR4_23(G4771,G4676,G4728,G2174,G1475);
  or OR4_24(G4772,G4729,G4730,G2175,G1476);
  or OR4_25(G4773,G4731,G4732,G2176,G1477);
  or OR4_26(G4774,G3055,G4509,G1497,G4747);
  and AND3_304(G4775,G4748,G1992,G2003);
  not NOT_784(G4776,G4681);
  not NOT_785(G4777,G4684);
  not NOT_786(G4778,G4687);
  and AND2_274(G4779,G4687,G1941);
  or OR3_42(G4780,G3087,G4750,G2340);
  or OR3_43(G4786,G3088,G4751,G2341);
  or OR3_44(G4792,G3089,G4752,G2342);
  or OR3_45(G4798,G3207,G4753,G2343);
  or OR3_46(G4804,G3091,G4754,G2345);
  or OR3_47(G4810,G3092,G4755,G2346);
  or OR3_48(G4816,G2887,G4756,G2347);
  or OR3_49(G4822,G3093,G4757,G2348);
  nand NAND2_325(G4828,G4761,G4691);
  nand NAND2_326(G4831,G4762,G4693);
  not NOT_787(G4834,G4694);
  nand NAND2_327(G4835,G4694,G4349);
  not NOT_788(G4836,G4697);
  nand NAND2_328(G4837,G4697,G4355);
  nand NAND2_329(G4838,G4763,G4701);
  nand NAND2_330(G4841,G4764,G4703);
  nand NAND2_331(G4844,G4765,G4705);
  not NOT_789(G4847,G4706);
  nand NAND2_332(G4848,G4706,G4374);
  and AND2_275(G4849,G4409,G4758);
  and AND2_276(G4850,G4758,G4606);
  and AND5_10(G4851,G156,G4776,G4777,G4264,G4377);
  and AND3_305(G4852,G4778,G1970,G1981);
  nand NAND2_333(G4853,G4125,G4834);
  nand NAND2_334(G4854,G4131,G4836);
  nand NAND2_335(G4855,G4170,G4847);
  and AND3_306(G4856,G4804,G1526,G1537);
  and AND3_307(G4857,G4780,G694,G1537);
  and AND3_308(G4858,G4810,G1526,G1537);
  and AND3_309(G4859,G4786,G694,G1537);
  and AND3_310(G4860,G4816,G1526,G1537);
  and AND3_311(G4861,G4792,G694,G1537);
  and AND3_312(G4862,G4822,G1526,G1537);
  and AND3_313(G4863,G4798,G694,G1537);
  and AND3_314(G4864,G4804,G1601,G1612);
  and AND3_315(G4865,G4780,G756,G1612);
  and AND3_316(G4866,G4810,G1601,G1612);
  and AND3_317(G4867,G4786,G756,G1612);
  and AND3_318(G4868,G4816,G1601,G1612);
  and AND3_319(G4869,G4792,G756,G1612);
  and AND3_320(G4870,G4822,G1601,G1612);
  and AND3_321(G4871,G4798,G756,G1612);
  and AND3_322(G4872,G4822,G1948,G1959);
  and AND3_323(G4873,G4798,G1218,G1959);
  and AND3_324(G4874,G4822,G1914,G1925);
  and AND3_325(G4875,G4798,G1184,G1925);
  and AND3_326(G4876,G4816,G1914,G1925);
  and AND3_327(G4877,G4792,G1184,G1925);
  and AND3_328(G4878,G4810,G1914,G1925);
  and AND3_329(G4879,G4786,G1184,G1925);
  and AND3_330(G4880,G4804,G1914,G1925);
  and AND3_331(G4881,G4780,G1184,G1925);
  and AND3_332(G4882,G4816,G1948,G1959);
  and AND3_333(G4883,G4792,G1218,G1959);
  and AND3_334(G4884,G4810,G1948,G1959);
  and AND3_335(G4885,G4786,G1218,G1959);
  and AND3_336(G4886,G4804,G1948,G1959);
  and AND3_337(G4887,G4780,G1218,G1959);
  not NOT_790(G4888,G4828);
  nand NAND2_336(G4889,G4828,G4230);
  not NOT_791(G4890,G4831);
  nand NAND2_337(G4891,G4831,G4233);
  nand NAND2_338(G4892,G4853,G4835);
  nand NAND2_339(G4895,G4854,G4837);
  not NOT_792(G4898,G4838);
  nand NAND2_340(G4899,G4838,G4244);
  not NOT_793(G4900,G4841);
  nand NAND2_341(G4901,G4841,G4246);
  not NOT_794(G4902,G4844);
  nand NAND2_342(G4903,G4844,G3694);
  nand NAND2_343(G4904,G4855,G4848);
  or OR4_27(G4907,G4856,G4857,G2158,G1461);
  or OR4_28(G4908,G4858,G4859,G2159,G1462);
  or OR4_29(G4909,G4860,G4861,G2160,G1463);
  or OR4_30(G4910,G4862,G4863,G2161,G1464);
  or OR4_31(G4911,G4864,G4865,G2169,G1470);
  or OR4_32(G4912,G4866,G4867,G2170,G1471);
  or OR4_33(G4913,G4868,G4869,G2171,G1472);
  or OR4_34(G4914,G4870,G4871,G2172,G1473);
  nand NAND2_344(G4915,G3939,G4888);
  nand NAND2_345(G4916,G3951,G4890);
  nand NAND2_346(G4917,G4008,G4898);
  nand NAND2_347(G4918,G4014,G4900);
  nand NAND2_348(G4919,G3256,G4902);
  nand NAND2_349(G4920,G4915,G4889);
  nand NAND2_350(G4923,G4916,G4891);
  not NOT_795(G4926,G4892);
  nand NAND2_351(G4927,G4892,G4236);
  not NOT_796(G4928,G4895);
  nand NAND2_352(G4929,G4895,G4241);
  nand NAND2_353(G4930,G4917,G4899);
  nand NAND2_354(G4933,G4918,G4901);
  nand NAND2_355(G4936,G4919,G4903);
  not NOT_797(G4939,G4904);
  nand NAND2_356(G4940,G4904,G3696);
  nand NAND2_357(G4941,G3963,G4926);
  nand NAND2_358(G4942,G3981,G4928);
  nand NAND2_359(G4943,G3262,G4939);
  not NOT_798(G4944,G4920);
  nand NAND2_360(G4945,G4920,G4231);
  not NOT_799(G4946,G4923);
  nand NAND2_361(G4947,G4923,G4234);
  nand NAND2_362(G4948,G4941,G4927);
  nand NAND2_363(G4951,G4942,G4929);
  not NOT_800(G4954,G4930);
  nand NAND2_364(G4955,G4930,G4245);
  not NOT_801(G4956,G4933);
  nand NAND2_365(G4957,G4933,G4247);
  not NOT_802(G4958,G4936);
  nand NAND2_366(G4959,G4936,G4248);
  nand NAND2_367(G4960,G4943,G4940);
  nand NAND2_368(G4963,G3942,G4944);
  nand NAND2_369(G4964,G3954,G4946);
  nand NAND2_370(G4965,G4011,G4954);
  nand NAND2_371(G4966,G4017,G4956);
  nand NAND2_372(G4967,G4020,G4958);
  nand NAND2_373(G4968,G4963,G4945);
  nand NAND2_374(G4971,G4964,G4947);
  not NOT_803(G4974,G4948);
  nand NAND2_375(G4975,G4948,G4237);
  not NOT_804(G4976,G4951);
  nand NAND2_376(G4977,G4951,G4242);
  nand NAND2_377(G4978,G4965,G4955);
  nand NAND2_378(G4981,G4966,G4957);
  nand NAND2_379(G4984,G4967,G4959);
  not NOT_805(G4987,G4960);
  nand NAND2_380(G4988,G4960,G4252);
  nand NAND2_381(G4989,G3966,G4974);
  nand NAND2_382(G4990,G3984,G4976);
  nand NAND2_383(G4991,G4029,G4987);
  not NOT_806(G4992,G4968);
  nand NAND2_384(G4993,G4968,G4232);
  not NOT_807(G4994,G4971);
  nand NAND2_385(G4995,G4971,G4235);
  nand NAND2_386(G4996,G4989,G4975);
  nand NAND2_387(G4999,G4990,G4977);
  not NOT_808(G5002,G4978);
  nand NAND2_388(G5003,G4978,G3691);
  not NOT_809(G5004,G4981);
  nand NAND2_389(G5005,G4981,G3693);
  not NOT_810(G5006,G4984);
  nand NAND2_390(G5007,G4984,G4249);
  nand NAND2_391(G5008,G4991,G4988);
  nand NAND2_392(G5011,G3945,G4992);
  nand NAND2_393(G5012,G3957,G4994);
  nand NAND2_394(G5013,G3241,G5002);
  nand NAND2_395(G5014,G3250,G5004);
  nand NAND2_396(G5015,G4023,G5006);
  nand NAND2_397(G5016,G5011,G4993);
  nand NAND2_398(G5019,G5012,G4995);
  not NOT_811(G5022,G4996);
  nand NAND2_399(G5023,G4996,G4238);
  not NOT_812(G5024,G4999);
  nand NAND2_400(G5025,G4999,G4243);
  nand NAND2_401(G5026,G5013,G5003);
  nand NAND2_402(G5029,G5014,G5005);
  nand NAND2_403(G5032,G5015,G5007);
  not NOT_813(G5035,G5008);
  nand NAND2_404(G5036,G5008,G4253);
  nand NAND2_405(G5037,G3969,G5022);
  nand NAND2_406(G5038,G3987,G5024);
  nand NAND2_407(G5039,G4032,G5035);
  not NOT_814(G5040,G5016);
  nand NAND2_408(G5041,G5016,G4200);
  not NOT_815(G5042,G5019);
  nand NAND2_409(G5043,G5019,G4201);
  not NOT_816(G5044,G5026);
  nand NAND2_410(G5045,G5026,G3664);
  not NOT_817(G5046,G5029);
  nand NAND2_411(G5047,G5029,G3665);
  nand NAND2_412(G5048,G5037,G5023);
  nand NAND2_413(G5051,G5038,G5025);
  not NOT_818(G5054,G5032);
  nand NAND2_414(G5055,G5032,G4250);
  nand NAND2_415(G5056,G5039,G5036);
  nand NAND2_416(G5059,G3948,G5040);
  nand NAND2_417(G5060,G3960,G5042);
  nand NAND2_418(G5061,G3244,G5044);
  nand NAND2_419(G5062,G3253,G5046);
  nand NAND2_420(G5063,G4026,G5054);
  nand NAND2_421(G5064,G5059,G5041);
  nand NAND2_422(G5067,G5060,G5043);
  nand NAND2_423(G5070,G5061,G5045);
  nand NAND2_424(G5073,G5062,G5047);
  not NOT_819(G5076,G5048);
  nand NAND2_425(G5077,G5048,G4239);
  not NOT_820(G5078,G5051);
  nand NAND2_426(G5079,G5051,G4240);
  nand NAND2_427(G5080,G5063,G5055);
  not NOT_821(G5083,G5056);
  nand NAND2_428(G5084,G5056,G4251);
  nand NAND2_429(G5085,G3972,G5076);
  nand NAND2_430(G5086,G3990,G5078);
  nand NAND2_431(G5087,G4035,G5083);
  and AND3_338(G5088,G5067,G4290,G690);
  and AND3_339(G5089,G5064,G4054,G690);
  and AND3_340(G5090,G5067,G4450,G157);
  and AND3_341(G5091,G5064,G4541,G157);
  not NOT_822(G5092,G5080);
  nand NAND2_432(G5093,G5080,G4075);
  and AND3_342(G5094,G5073,G4316,G752);
  and AND3_343(G5095,G5070,G4068,G752);
  and AND3_344(G5096,G5073,G4473,G162);
  and AND3_345(G5097,G5070,G4546,G162);
  nand NAND2_433(G5098,G5085,G5077);
  nand NAND2_434(G5101,G5086,G5079);
  nand NAND2_435(G5104,G5087,G5084);
  nand NAND2_436(G5107,G3745,G5092);
  or OR4_35(G5108,G5088,G5089,G5090,G5091);
  or OR4_36(G5111,G5094,G5095,G5096,G5097);
  not NOT_823(G5114,G5098);
  nand NAND2_437(G5115,G5098,G4202);
  not NOT_824(G5116,G5101);
  nand NAND2_438(G5117,G5101,G4203);
  nand NAND2_439(G5118,G5107,G5093);
  not NOT_825(G5119,G5104);
  nand NAND2_440(G5120,G5104,G4076);
  nand NAND2_441(G5121,G3975,G5114);
  nand NAND2_442(G5122,G3978,G5116);
  not NOT_826(G5123,G5108);
  nand NAND2_443(G5124,G3748,G5119);
  and AND2_277(G5125,G162,G5118);
  not NOT_827(G5126,G5111);
  nand NAND2_444(G5127,G5121,G5115);
  nand NAND2_445(G5128,G5122,G5117);
  nand NAND2_446(G5129,G5124,G5120);
  not NOT_828(G5130,G5128);
  and AND2_278(G5131,G157,G5127);
  not NOT_829(G5132,G5129);
  and AND2_279(G5133,G5130,G690);
  and AND2_280(G5134,G5132,G752);
  or OR2_82(G5135,G5133,G5131);
  or OR2_83(G5138,G5134,G5125);
  nand NAND2_447(G5141,G5135,G5123);
  not NOT_830(G5142,G5135);
  nand NAND2_448(G5143,G5138,G5126);
  not NOT_831(G5144,G5138);
  nand NAND2_449(G5145,G5108,G5142);
  nand NAND2_450(G5146,G5111,G5144);
  nand NAND2_451(G5147,G5141,G5145);
  nand NAND2_452(G5150,G5143,G5146);
  and AND3_346(G5153,G5150,G1264,G2003);
  and AND3_347(G5154,G5147,G1248,G1981);
  not NOT_832(G5155,G5147);
  not NOT_833(G5156,G5150);
  and AND2_281(G5157,G5155,G1214);
  and AND2_282(G5158,G5156,G1214);
  or OR2_84(G5159,G4779,G5157);
  or OR2_85(G5162,G4749,G5158);
  and AND2_283(G5165,G5159,G1936);
  and AND2_284(G5166,G5162,G1936);
  and AND2_285(G5167,G5159,G1936);
  and AND2_286(G5168,G5162,G1936);
  or OR2_86(G5169,G5165,G1944);
  or OR2_87(G5172,G5166,G1945);
  or OR2_88(G5175,G5167,G1946);
  or OR2_89(G5178,G5168,G1947);
  and AND3_348(G5181,G5178,G1652,G1663);
  and AND3_349(G5182,G5175,G860,G1663);
  and AND3_350(G5183,G5178,G1674,G1685);
  and AND3_351(G5184,G5175,G884,G1685);
  and AND3_352(G5185,G5172,G1554,G1565);
  and AND3_353(G5186,G5169,G718,G1565);
  and AND3_354(G5187,G5172,G1629,G1640);
  and AND3_355(G5188,G5169,G780,G1640);
  or OR4_37(G5189,G5185,G5186,G2203,G1576);
  or OR4_38(G5190,G5187,G5188,G2204,G1651);
  and AND2_287(G5191,G5189,G1548);
  and AND2_288(G5192,G5190,G1623);
  not NOT_834(G5193,G66);
  not NOT_835(G5194,G113);
  not NOT_836(G5195,G165);
  not NOT_837(G5196,G151);
  not NOT_838(G5197,G127);
  not NOT_839(G5198,G131);
  and AND2_289(G5199,G153,G156);
  not NOT_840(G5200,G152);
  not NOT_841(G5201,G151);
  not NOT_842(G5202,G151);
  not NOT_843(G5203,G125);
  not NOT_844(G5204,G129);
  and AND2_290(G5205,G66,G67);
  not NOT_845(G5206,G99);
  not NOT_846(G5207,G153);
  not NOT_847(G5208,G156);
  not NOT_848(G5209,G155);
  not NOT_849(G5210,G684);
  and AND2_291(G5211,G63,G685);
  not NOT_850(G5212,G687);
  not NOT_851(G5213,G688);
  not NOT_852(G5214,G742);
  not NOT_853(G5215,G749);
  not NOT_854(G5216,G980);
  not NOT_855(G5217,G1067);
  not NOT_856(G5218,G1308);
  not NOT_857(G5219,G1067);
  nand NAND2_453(G5220,G976,G65);
  not NOT_858(G5221,G976);
  not NOT_859(G5222,G1577);
  not NOT_860(G5223,G1577);
  not NOT_861(G5224,G1577);
  not NOT_862(G5225,G1577);
  not NOT_863(G5226,G2064);
  not NOT_864(G5227,G2064);
  not NOT_865(G5228,G2528);
  not NOT_866(G5229,G2533);
  not NOT_867(G5230,G2538);
  not NOT_868(G5231,G2539);
  and AND2_292(G5232,G2671,G1750);
  and AND2_293(G5233,G2672,G1750);
  and AND2_294(G5234,G2673,G1750);
  and AND2_295(G5235,G2674,G1750);
  and AND3_356(G5236,G3105,G3106,G2669);
  and AND3_357(G5237,G3107,G3108,G3281);
  and AND2_296(G5238,G3793,G3802);
  and AND2_297(G5239,G3825,G3834);
  and AND2_298(G5240,G3852,G3859);
  and AND2_299(G5241,G3765,G3776);
  not NOT_869(G5242,G4077);
  not NOT_870(G5243,G4227);
  or OR2_90(G5244,G4044,G4260);
  or OR2_91(G5245,G4045,G4261);
  or OR2_92(G5246,G4046,G4262);
  or OR2_93(G5247,G4047,G4263);
  not NOT_871(G5248,G4323);
  not NOT_872(G5249,G4562);
  not NOT_873(G5250,G4554);
  not NOT_874(G5251,G4606);
  or OR4_39(G5252,G4425,G4677,G2182,G1479);
  not NOT_875(G5253,G4664);
  not NOT_876(G5254,G4648);
  not NOT_877(G5255,G4642);
  or OR4_40(G5256,G4426,G4680,G2201,G1499);
  not NOT_878(G5257,G4658);
  not NOT_879(G5258,G4636);
  not NOT_880(G5259,G4630);
  not NOT_881(G5260,G4624);
  not NOT_882(G5261,G4681);
  not NOT_883(G5262,G4684);
  and AND9_0(G5263,G4507,G4530,G4531,G4532,G4533,G4709,G4710,G4711,G4712);
  and AND9_1(G5264,G4183,G4508,G4534,G4535,G4536,G4713,G4714,G4715,G4716);
  and AND2_300(G5265,G4719,G1548);
  and AND2_301(G5266,G4727,G1623);
  or OR4_41(G5267,G4733,G4734,G2187,G1484);
  or OR4_42(G5268,G4735,G4736,G2188,G1485);
  or OR4_43(G5269,G4737,G4738,G2189,G1486);
  or OR4_44(G5270,G4678,G4739,G2190,G1487);
  or OR4_45(G5271,G4740,G4741,G2195,G1492);
  or OR4_46(G5272,G4742,G4743,G2196,G1493);
  or OR4_47(G5273,G4744,G4745,G2197,G1494);
  or OR4_48(G5274,G4679,G4746,G2198,G1495);
  and AND2_302(G5275,G4766,G1520);
  and AND2_303(G5276,G4767,G1548);
  and AND2_304(G5277,G4768,G1548);
  and AND2_305(G5278,G4769,G1548);
  and AND2_306(G5279,G4770,G1595);
  and AND2_307(G5280,G4771,G1623);
  and AND2_308(G5281,G4772,G1623);
  and AND2_309(G5282,G4773,G1623);
  and AND2_310(G5283,G686,G4774);
  or OR2_94(G5284,G4849,G4850);
  not NOT_884(G5285,G4822);
  not NOT_885(G5286,G4816);
  not NOT_886(G5287,G4810);
  not NOT_887(G5288,G4804);
  and AND3_358(G5289,G689,G4851,G99);
  not NOT_888(G5290,G4798);
  not NOT_889(G5291,G4792);
  not NOT_890(G5292,G4786);
  not NOT_891(G5293,G4780);
  or OR4_49(G5294,G4872,G4873,G2179,G1478);
  or OR4_50(G5295,G4874,G4875,G2183,G1480);
  or OR4_51(G5296,G4876,G4877,G2184,G1481);
  or OR4_52(G5297,G4878,G4879,G2185,G1482);
  or OR4_53(G5298,G4880,G4881,G2186,G1483);
  or OR4_54(G5299,G4882,G4883,G2192,G1489);
  or OR4_55(G5300,G4884,G4885,G2193,G1490);
  or OR4_56(G5301,G4886,G4887,G2194,G1491);
  and AND2_311(G5302,G4907,G1520);
  and AND2_312(G5303,G4908,G1520);
  and AND2_313(G5304,G4909,G1520);
  and AND2_314(G5305,G4910,G1520);
  and AND2_315(G5306,G4911,G1595);
  and AND2_316(G5307,G4912,G1595);
  and AND2_317(G5308,G4913,G1595);
  and AND2_318(G5309,G4914,G1595);
  or OR4_57(G5310,G4775,G5153,G2200,G1498);
  or OR4_58(G5311,G4852,G5154,G2202,G1500);
  or OR4_59(G5312,G5181,G5182,G2191,G1488);
  or OR4_60(G5313,G5183,G5184,G2199,G1496);
  not NOT_892(G5314,G5191);
  not NOT_893(G5315,G5192);

endmodule

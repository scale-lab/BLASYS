module sin_tb;
reg [23:0] pi;
wire [24:0] po;
sin dut(pi[0], pi[1], pi[2], pi[3], pi[4], pi[5], pi[6], pi[7], pi[8], pi[9], pi[10], pi[11], pi[12], pi[13], pi[14], pi[15], pi[16], pi[17], pi[18], pi[19], pi[20], pi[21], pi[22], pi[23], po[0], po[1], po[2], po[3], po[4], po[5], po[6], po[7], po[8], po[9], po[10], po[11], po[12], po[13], po[14], po[15], po[16], po[17], po[18], po[19], po[20], po[21], po[22], po[23], po[24]);
initial
begin
# 1  pi=24'b101011000010101111111011;
#1 $display("%b", po);
# 1  pi=24'b000101100010000011110100;
#1 $display("%b", po);
# 1  pi=24'b001011001001110001101111;
#1 $display("%b", po);
# 1  pi=24'b101100100010110111000001;
#1 $display("%b", po);
# 1  pi=24'b110110001101100111000100;
#1 $display("%b", po);
# 1  pi=24'b100010110011110110110110;
#1 $display("%b", po);
# 1  pi=24'b000111111101000011000111;
#1 $display("%b", po);
# 1  pi=24'b010100011000100100111000;
#1 $display("%b", po);
# 1  pi=24'b100110011100000000100000;
#1 $display("%b", po);
# 1  pi=24'b110110001000001011110111;
#1 $display("%b", po);
# 1  pi=24'b100010100110100011101110;
#1 $display("%b", po);
# 1  pi=24'b100100000111101101010101;
#1 $display("%b", po);
# 1  pi=24'b011010100100111111111001;
#1 $display("%b", po);
# 1  pi=24'b010111001000001111011010;
#1 $display("%b", po);
# 1  pi=24'b000010011010110000110110;
#1 $display("%b", po);
# 1  pi=24'b110000000100011101100001;
#1 $display("%b", po);
# 1  pi=24'b101001100011010001101100;
#1 $display("%b", po);
# 1  pi=24'b010010001101111010011110;
#1 $display("%b", po);
# 1  pi=24'b111011111100111101010100;
#1 $display("%b", po);
# 1  pi=24'b111101110000100011001001;
#1 $display("%b", po);
# 1  pi=24'b111110101011000100101110;
#1 $display("%b", po);
# 1  pi=24'b110001010010110100001001;
#1 $display("%b", po);
# 1  pi=24'b101111000110011101011011;
#1 $display("%b", po);
# 1  pi=24'b000000001111000100110010;
#1 $display("%b", po);
# 1  pi=24'b010011110101011110000010;
#1 $display("%b", po);
# 1  pi=24'b110111001010100001010010;
#1 $display("%b", po);
# 1  pi=24'b111100110110110011001100;
#1 $display("%b", po);
# 1  pi=24'b110010011111010111010001;
#1 $display("%b", po);
# 1  pi=24'b000111111010011111001001;
#1 $display("%b", po);
# 1  pi=24'b000010101110110001011110;
#1 $display("%b", po);
# 1  pi=24'b010001010100010010100101;
#1 $display("%b", po);
# 1  pi=24'b011100110001000001010000;
#1 $display("%b", po);
# 1  pi=24'b011101100110011001000011;
#1 $display("%b", po);
# 1  pi=24'b101101110000100100100111;
#1 $display("%b", po);
# 1  pi=24'b111001100100100011000101;
#1 $display("%b", po);
# 1  pi=24'b001111000000000010110000;
#1 $display("%b", po);
# 1  pi=24'b100110110100100011111111;
#1 $display("%b", po);
# 1  pi=24'b101111010001011000001010;
#1 $display("%b", po);
# 1  pi=24'b110111010100110000111101;
#1 $display("%b", po);
# 1  pi=24'b000011101010001001001110;
#1 $display("%b", po);
# 1  pi=24'b011010111001010010100110;
#1 $display("%b", po);
# 1  pi=24'b000010101010110110001110;
#1 $display("%b", po);
# 1  pi=24'b001001101011000101111101;
#1 $display("%b", po);
# 1  pi=24'b110001001100001111000110;
#1 $display("%b", po);
# 1  pi=24'b110000011011000010101010;
#1 $display("%b", po);
# 1  pi=24'b010011010100110110011100;
#1 $display("%b", po);
# 1  pi=24'b110001010000010001011000;
#1 $display("%b", po);
# 1  pi=24'b100010000011000011110100;
#1 $display("%b", po);
# 1  pi=24'b001101001010111011010111;
#1 $display("%b", po);
# 1  pi=24'b111010000001110110100001;
#1 $display("%b", po);
# 1  pi=24'b001110011100100110010111;
#1 $display("%b", po);
# 1  pi=24'b111011001100101011110000;
#1 $display("%b", po);
# 1  pi=24'b011010100001000010011100;
#1 $display("%b", po);
# 1  pi=24'b001001111110001101011100;
#1 $display("%b", po);
# 1  pi=24'b101000010011001110010001;
#1 $display("%b", po);
# 1  pi=24'b101101001001111100100000;
#1 $display("%b", po);
# 1  pi=24'b011010100010101001000111;
#1 $display("%b", po);
# 1  pi=24'b001001011011101101110011;
#1 $display("%b", po);
# 1  pi=24'b011000001101100111010010;
#1 $display("%b", po);
# 1  pi=24'b101000110001001100111100;
#1 $display("%b", po);
# 1  pi=24'b000010000100010010101101;
#1 $display("%b", po);
# 1  pi=24'b000111111111011010100100;
#1 $display("%b", po);
# 1  pi=24'b010101101000100001101100;
#1 $display("%b", po);
# 1  pi=24'b001100010011101111011010;
#1 $display("%b", po);
# 1  pi=24'b110011011101111001000011;
#1 $display("%b", po);
# 1  pi=24'b110010101001010010111101;
#1 $display("%b", po);
# 1  pi=24'b010000111011110011111110;
#1 $display("%b", po);
# 1  pi=24'b011100010101101010011100;
#1 $display("%b", po);
# 1  pi=24'b011010011100111110110101;
#1 $display("%b", po);
# 1  pi=24'b101000001001100101111010;
#1 $display("%b", po);
# 1  pi=24'b100110100101000101011101;
#1 $display("%b", po);
# 1  pi=24'b100101011110001100101000;
#1 $display("%b", po);
# 1  pi=24'b101011010111001000100100;
#1 $display("%b", po);
# 1  pi=24'b000110011000000010001111;
#1 $display("%b", po);
# 1  pi=24'b011000010011111000001001;
#1 $display("%b", po);
# 1  pi=24'b010111011000010100110010;
#1 $display("%b", po);
# 1  pi=24'b110110100110110000010000;
#1 $display("%b", po);
# 1  pi=24'b101011000001001000010010;
#1 $display("%b", po);
# 1  pi=24'b011100110000100100111110;
#1 $display("%b", po);
# 1  pi=24'b001111011010001011010011;
#1 $display("%b", po);
# 1  pi=24'b111110001111101010001100;
#1 $display("%b", po);
# 1  pi=24'b001000111011100010011111;
#1 $display("%b", po);
# 1  pi=24'b100010100001111011111100;
#1 $display("%b", po);
# 1  pi=24'b010001111101110111101011;
#1 $display("%b", po);
# 1  pi=24'b101010010010100011001100;
#1 $display("%b", po);
# 1  pi=24'b001101110001111110011011;
#1 $display("%b", po);
# 1  pi=24'b011110101110111001011110;
#1 $display("%b", po);
# 1  pi=24'b100001101100010010110101;
#1 $display("%b", po);
# 1  pi=24'b000101111001011100101111;
#1 $display("%b", po);
# 1  pi=24'b001000101111010111011100;
#1 $display("%b", po);
# 1  pi=24'b101000110101010110010101;
#1 $display("%b", po);
# 1  pi=24'b010010111110111011100111;
#1 $display("%b", po);
# 1  pi=24'b101100001011110000001101;
#1 $display("%b", po);
# 1  pi=24'b001000000101010001100000;
#1 $display("%b", po);
# 1  pi=24'b010101011001111100010001;
#1 $display("%b", po);
# 1  pi=24'b100110101101010110100001;
#1 $display("%b", po);
# 1  pi=24'b010110000101111001001110;
#1 $display("%b", po);
# 1  pi=24'b100011011001101000111000;
#1 $display("%b", po);
# 1  pi=24'b111100001011001110001001;
#1 $display("%b", po);
# 1  pi=24'b001101001100101011010111;
#1 $display("%b", po);
# 1  pi=24'b000001101100000111100101;
#1 $display("%b", po);
# 1  pi=24'b101011001000011110101101;
#1 $display("%b", po);
# 1  pi=24'b010010010001010010010101;
#1 $display("%b", po);
# 1  pi=24'b101010011110110110110100;
#1 $display("%b", po);
# 1  pi=24'b000011010101101110100110;
#1 $display("%b", po);
# 1  pi=24'b101011000111001110011001;
#1 $display("%b", po);
# 1  pi=24'b011111000010101011011001;
#1 $display("%b", po);
# 1  pi=24'b101011010011101111111001;
#1 $display("%b", po);
# 1  pi=24'b010110110111110001001001;
#1 $display("%b", po);
# 1  pi=24'b111001101101000101111001;
#1 $display("%b", po);
# 1  pi=24'b011111100100100011011110;
#1 $display("%b", po);
# 1  pi=24'b110101110101110110111000;
#1 $display("%b", po);
# 1  pi=24'b100010011101100010101100;
#1 $display("%b", po);
# 1  pi=24'b001010011111010101111010;
#1 $display("%b", po);
# 1  pi=24'b100100111000010001010101;
#1 $display("%b", po);
# 1  pi=24'b011010110101110100010000;
#1 $display("%b", po);
# 1  pi=24'b101101011110010111111100;
#1 $display("%b", po);
# 1  pi=24'b011010100001110100101101;
#1 $display("%b", po);
# 1  pi=24'b000001110010110101110001;
#1 $display("%b", po);
# 1  pi=24'b100010001110001000111000;
#1 $display("%b", po);
# 1  pi=24'b001101110010110111110100;
#1 $display("%b", po);
# 1  pi=24'b100110011110100100100001;
#1 $display("%b", po);
# 1  pi=24'b000100110111000101110101;
#1 $display("%b", po);
# 1  pi=24'b111110000110001001011011;
#1 $display("%b", po);
# 1  pi=24'b100100100101000011000100;
#1 $display("%b", po);
# 1  pi=24'b001110000000001001000101;
#1 $display("%b", po);
# 1  pi=24'b101100101010101111111110;
#1 $display("%b", po);
# 1  pi=24'b010111000000100000011010;
#1 $display("%b", po);
# 1  pi=24'b100110101100000110110011;
#1 $display("%b", po);
# 1  pi=24'b011000001101101100101000;
#1 $display("%b", po);
# 1  pi=24'b000000000000111110110010;
#1 $display("%b", po);
# 1  pi=24'b111011011000011000010110;
#1 $display("%b", po);
# 1  pi=24'b100100110111111000100001;
#1 $display("%b", po);
# 1  pi=24'b000010101011000100110001;
#1 $display("%b", po);
# 1  pi=24'b000101100100101011101010;
#1 $display("%b", po);
# 1  pi=24'b111010000100101101111010;
#1 $display("%b", po);
# 1  pi=24'b111000110000000100111110;
#1 $display("%b", po);
# 1  pi=24'b011101110101110011101100;
#1 $display("%b", po);
# 1  pi=24'b101001100100110100001001;
#1 $display("%b", po);
# 1  pi=24'b001010010011111111111111;
#1 $display("%b", po);
# 1  pi=24'b010101011100111101100011;
#1 $display("%b", po);
# 1  pi=24'b011111011100000000000110;
#1 $display("%b", po);
# 1  pi=24'b000111011010011110101001;
#1 $display("%b", po);
# 1  pi=24'b010000010101101010110001;
#1 $display("%b", po);
# 1  pi=24'b111011100011110011100100;
#1 $display("%b", po);
# 1  pi=24'b100010111111000101100101;
#1 $display("%b", po);
# 1  pi=24'b100101101010110111000001;
#1 $display("%b", po);
# 1  pi=24'b101101111110110111101110;
#1 $display("%b", po);
# 1  pi=24'b011010110000001001011100;
#1 $display("%b", po);
# 1  pi=24'b010011001001101100100100;
#1 $display("%b", po);
# 1  pi=24'b010000001010001101100101;
#1 $display("%b", po);
# 1  pi=24'b101001011110010001101100;
#1 $display("%b", po);
# 1  pi=24'b010011100001110100011011;
#1 $display("%b", po);
# 1  pi=24'b000010001111100010011111;
#1 $display("%b", po);
# 1  pi=24'b101011110001010011100010;
#1 $display("%b", po);
# 1  pi=24'b000111100011011110101010;
#1 $display("%b", po);
# 1  pi=24'b011101011000001110101101;
#1 $display("%b", po);
# 1  pi=24'b011100001111100011101001;
#1 $display("%b", po);
# 1  pi=24'b000110110010010111011010;
#1 $display("%b", po);
# 1  pi=24'b101101101111110000100010;
#1 $display("%b", po);
# 1  pi=24'b101100110101101101111101;
#1 $display("%b", po);
# 1  pi=24'b101110111010010101000101;
#1 $display("%b", po);
# 1  pi=24'b010100100000001010011100;
#1 $display("%b", po);
# 1  pi=24'b001101000101011110101010;
#1 $display("%b", po);
# 1  pi=24'b111011000001111010101110;
#1 $display("%b", po);
# 1  pi=24'b101010001111011100101011;
#1 $display("%b", po);
# 1  pi=24'b101111110010100111110101;
#1 $display("%b", po);
# 1  pi=24'b111111000101110100101111;
#1 $display("%b", po);
# 1  pi=24'b101011000001011101110101;
#1 $display("%b", po);
# 1  pi=24'b101000101011001101010010;
#1 $display("%b", po);
# 1  pi=24'b111001001110111110110111;
#1 $display("%b", po);
# 1  pi=24'b011011010111100110111110;
#1 $display("%b", po);
# 1  pi=24'b110111110000011010001010;
#1 $display("%b", po);
# 1  pi=24'b110000101111000010010110;
#1 $display("%b", po);
# 1  pi=24'b101001111111110001101100;
#1 $display("%b", po);
# 1  pi=24'b101110111100010110000111;
#1 $display("%b", po);
# 1  pi=24'b110110010110110001100111;
#1 $display("%b", po);
# 1  pi=24'b100110000100000101111110;
#1 $display("%b", po);
# 1  pi=24'b111010110011101100011011;
#1 $display("%b", po);
# 1  pi=24'b100110011010101000000010;
#1 $display("%b", po);
# 1  pi=24'b010000111001010011011110;
#1 $display("%b", po);
# 1  pi=24'b100010011010001101000100;
#1 $display("%b", po);
# 1  pi=24'b101110100001001111110111;
#1 $display("%b", po);
# 1  pi=24'b011010001001000011001001;
#1 $display("%b", po);
# 1  pi=24'b001111110000011111110010;
#1 $display("%b", po);
# 1  pi=24'b000101000111010000100100;
#1 $display("%b", po);
# 1  pi=24'b111000011111101011101110;
#1 $display("%b", po);
# 1  pi=24'b001000000000110111100101;
#1 $display("%b", po);
# 1  pi=24'b100111000011010101001000;
#1 $display("%b", po);
# 1  pi=24'b000001111100001100100110;
#1 $display("%b", po);
# 1  pi=24'b100000000010011010100011;
#1 $display("%b", po);
# 1  pi=24'b110111110111111011100000;
#1 $display("%b", po);
# 1  pi=24'b001000011100000001100000;
#1 $display("%b", po);
# 1  pi=24'b100001111001001010011100;
#1 $display("%b", po);
# 1  pi=24'b100011111101010011000010;
#1 $display("%b", po);
# 1  pi=24'b101100110011010011111101;
#1 $display("%b", po);
# 1  pi=24'b111011001000001111000100;
#1 $display("%b", po);
# 1  pi=24'b110111001111000111100100;
#1 $display("%b", po);
# 1  pi=24'b001111110000110100001111;
#1 $display("%b", po);
# 1  pi=24'b110111001111111100110010;
#1 $display("%b", po);
# 1  pi=24'b110100101101010011101011;
#1 $display("%b", po);
# 1  pi=24'b101111010011011010011111;
#1 $display("%b", po);
# 1  pi=24'b010010001101001001000100;
#1 $display("%b", po);
# 1  pi=24'b101100111100001111000111;
#1 $display("%b", po);
# 1  pi=24'b110011101110001000111110;
#1 $display("%b", po);
# 1  pi=24'b100110101101011111100100;
#1 $display("%b", po);
# 1  pi=24'b101001011000101001011100;
#1 $display("%b", po);
# 1  pi=24'b101011110001000011000011;
#1 $display("%b", po);
# 1  pi=24'b010010100010100011100101;
#1 $display("%b", po);
# 1  pi=24'b111011001001001010101010;
#1 $display("%b", po);
# 1  pi=24'b100101100000010001011110;
#1 $display("%b", po);
# 1  pi=24'b110100111010001111110011;
#1 $display("%b", po);
# 1  pi=24'b011011010110010001111010;
#1 $display("%b", po);
# 1  pi=24'b000101110110001000010111;
#1 $display("%b", po);
# 1  pi=24'b111101100100010000100001;
#1 $display("%b", po);
# 1  pi=24'b110100011110000010011011;
#1 $display("%b", po);
# 1  pi=24'b010101111011011110001001;
#1 $display("%b", po);
# 1  pi=24'b101010000010010010111100;
#1 $display("%b", po);
# 1  pi=24'b100010100100010010010000;
#1 $display("%b", po);
# 1  pi=24'b100100000111110001001001;
#1 $display("%b", po);
# 1  pi=24'b010000101100111100011100;
#1 $display("%b", po);
# 1  pi=24'b010010010111111111001000;
#1 $display("%b", po);
# 1  pi=24'b101010011110000001011000;
#1 $display("%b", po);
# 1  pi=24'b000101110100100000111111;
#1 $display("%b", po);
# 1  pi=24'b111010011110001101101111;
#1 $display("%b", po);
# 1  pi=24'b000001101010111011000010;
#1 $display("%b", po);
# 1  pi=24'b011101001110111100010001;
#1 $display("%b", po);
# 1  pi=24'b010000011000100101000110;
#1 $display("%b", po);
# 1  pi=24'b110000101101000111000000;
#1 $display("%b", po);
# 1  pi=24'b101110011010011010000110;
#1 $display("%b", po);
# 1  pi=24'b111010111010011100000101;
#1 $display("%b", po);
# 1  pi=24'b010001101011011100101101;
#1 $display("%b", po);
# 1  pi=24'b011000100010001111101011;
#1 $display("%b", po);
# 1  pi=24'b100110101101011001010110;
#1 $display("%b", po);
# 1  pi=24'b011000110100010000110100;
#1 $display("%b", po);
# 1  pi=24'b100110100000001110000011;
#1 $display("%b", po);
# 1  pi=24'b010111001011010010100110;
#1 $display("%b", po);
# 1  pi=24'b100010010011011111010100;
#1 $display("%b", po);
# 1  pi=24'b010010010000101100111100;
#1 $display("%b", po);
# 1  pi=24'b101011101010010010011001;
#1 $display("%b", po);
# 1  pi=24'b101011010011101001011000;
#1 $display("%b", po);
# 1  pi=24'b010010001011000100111100;
#1 $display("%b", po);
# 1  pi=24'b100000110001000000000110;
#1 $display("%b", po);
# 1  pi=24'b101101001011110111101010;
#1 $display("%b", po);
# 1  pi=24'b100011110000101101111111;
#1 $display("%b", po);
# 1  pi=24'b101100000011111111010110;
#1 $display("%b", po);
# 1  pi=24'b001000100010101101000100;
#1 $display("%b", po);
# 1  pi=24'b111001000111011000110110;
#1 $display("%b", po);
# 1  pi=24'b011010000100000010101010;
#1 $display("%b", po);
# 1  pi=24'b111101010100110100110110;
#1 $display("%b", po);
# 1  pi=24'b000100111011000100010100;
#1 $display("%b", po);
# 1  pi=24'b111100100111101111001110;
#1 $display("%b", po);
# 1  pi=24'b011001011110010011000001;
#1 $display("%b", po);
# 1  pi=24'b101010101000010110011000;
#1 $display("%b", po);
# 1  pi=24'b100001001101101011010010;
#1 $display("%b", po);
# 1  pi=24'b010111101011011001010110;
#1 $display("%b", po);
# 1  pi=24'b100011000001010100000100;
#1 $display("%b", po);
# 1  pi=24'b100011000010010011111010;
#1 $display("%b", po);
# 1  pi=24'b110000011100011100001101;
#1 $display("%b", po);
# 1  pi=24'b110011010011000101100101;
#1 $display("%b", po);
# 1  pi=24'b000101001000111111100101;
#1 $display("%b", po);
# 1  pi=24'b111010100001101101101101;
#1 $display("%b", po);
# 1  pi=24'b010000011011010100100101;
#1 $display("%b", po);
# 1  pi=24'b100011011110001101011011;
#1 $display("%b", po);
# 1  pi=24'b100000010011101000001101;
#1 $display("%b", po);
# 1  pi=24'b100010010111011100110011;
#1 $display("%b", po);
# 1  pi=24'b000111001010111100110111;
#1 $display("%b", po);
# 1  pi=24'b101111001001110010010010;
#1 $display("%b", po);
# 1  pi=24'b011011101011100101111111;
#1 $display("%b", po);
# 1  pi=24'b111111001101011010110111;
#1 $display("%b", po);
# 1  pi=24'b011001110101001100100111;
#1 $display("%b", po);
# 1  pi=24'b010100000001001110101000;
#1 $display("%b", po);
# 1  pi=24'b001111100000100001001100;
#1 $display("%b", po);
# 1  pi=24'b101010101001000001110111;
#1 $display("%b", po);
# 1  pi=24'b110001111101101100001001;
#1 $display("%b", po);
# 1  pi=24'b111111010001010010011001;
#1 $display("%b", po);
# 1  pi=24'b000010011010100110101101;
#1 $display("%b", po);
# 1  pi=24'b010010001001100010010010;
#1 $display("%b", po);
# 1  pi=24'b110100000010001101101010;
#1 $display("%b", po);
# 1  pi=24'b010111011111001111111010;
#1 $display("%b", po);
# 1  pi=24'b100100100100111000000000;
#1 $display("%b", po);
# 1  pi=24'b010100111110110111000001;
#1 $display("%b", po);
# 1  pi=24'b010010100011100101110001;
#1 $display("%b", po);
# 1  pi=24'b010001001000101000100101;
#1 $display("%b", po);
# 1  pi=24'b011001111011011000011110;
#1 $display("%b", po);
# 1  pi=24'b010011111010101011100110;
#1 $display("%b", po);
# 1  pi=24'b111000010101101110110111;
#1 $display("%b", po);
# 1  pi=24'b011111111010001100010110;
#1 $display("%b", po);
# 1  pi=24'b001111011110110111101011;
#1 $display("%b", po);
# 1  pi=24'b101111001111000001000110;
#1 $display("%b", po);
# 1  pi=24'b011011100110101100001111;
#1 $display("%b", po);
# 1  pi=24'b101111010011000101000011;
#1 $display("%b", po);
# 1  pi=24'b001110010110000100100010;
#1 $display("%b", po);
# 1  pi=24'b110001011000011001101011;
#1 $display("%b", po);
# 1  pi=24'b001000100000010010010001;
#1 $display("%b", po);
# 1  pi=24'b000001100110000000010011;
#1 $display("%b", po);
# 1  pi=24'b111111011100100000111101;
#1 $display("%b", po);
# 1  pi=24'b011000101000000000000101;
#1 $display("%b", po);
# 1  pi=24'b001100011100110100011000;
#1 $display("%b", po);
# 1  pi=24'b100111011111101000101110;
#1 $display("%b", po);
# 1  pi=24'b111101001111110011010000;
#1 $display("%b", po);
# 1  pi=24'b110010011111000111010100;
#1 $display("%b", po);
# 1  pi=24'b111001110011000001111100;
#1 $display("%b", po);
# 1  pi=24'b100011100100110110000011;
#1 $display("%b", po);
# 1  pi=24'b101100110000110010000011;
#1 $display("%b", po);
# 1  pi=24'b010000100101100001101111;
#1 $display("%b", po);
# 1  pi=24'b000010101001100010111000;
#1 $display("%b", po);
# 1  pi=24'b101111111111101001100100;
#1 $display("%b", po);
# 1  pi=24'b001111100010100000000101;
#1 $display("%b", po);
# 1  pi=24'b101111010001010011001110;
#1 $display("%b", po);
# 1  pi=24'b010111111110010001111010;
#1 $display("%b", po);
# 1  pi=24'b010010111001101111101100;
#1 $display("%b", po);
# 1  pi=24'b101010111101001101111110;
#1 $display("%b", po);
# 1  pi=24'b100001001100100010110010;
#1 $display("%b", po);
# 1  pi=24'b001000011110000110101101;
#1 $display("%b", po);
# 1  pi=24'b111100001110101011110000;
#1 $display("%b", po);
# 1  pi=24'b011000001001111110110110;
#1 $display("%b", po);
# 1  pi=24'b100100101101111010000100;
#1 $display("%b", po);
# 1  pi=24'b001011001100000010101000;
#1 $display("%b", po);
# 1  pi=24'b000011111001001010110111;
#1 $display("%b", po);
# 1  pi=24'b001011001010010100000000;
#1 $display("%b", po);
# 1  pi=24'b000011100100010001011000;
#1 $display("%b", po);
# 1  pi=24'b001010000110111100100000;
#1 $display("%b", po);
# 1  pi=24'b001011111111000111011101;
#1 $display("%b", po);
# 1  pi=24'b100110111100101100110101;
#1 $display("%b", po);
# 1  pi=24'b000001001100110101000110;
#1 $display("%b", po);
# 1  pi=24'b000000001100111001100001;
#1 $display("%b", po);
# 1  pi=24'b011111110100011001101010;
#1 $display("%b", po);
# 1  pi=24'b010011001001101011010000;
#1 $display("%b", po);
# 1  pi=24'b101101011011110001010001;
#1 $display("%b", po);
# 1  pi=24'b111010001000000000010001;
#1 $display("%b", po);
# 1  pi=24'b011110010001001101100010;
#1 $display("%b", po);
# 1  pi=24'b001011000110100101000111;
#1 $display("%b", po);
# 1  pi=24'b100110011111000010011000;
#1 $display("%b", po);
# 1  pi=24'b001011000010001010010110;
#1 $display("%b", po);
# 1  pi=24'b000100001101011000001011;
#1 $display("%b", po);
# 1  pi=24'b010000010111011110111111;
#1 $display("%b", po);
# 1  pi=24'b000111101001111011111111;
#1 $display("%b", po);
# 1  pi=24'b001010110000001011101110;
#1 $display("%b", po);
# 1  pi=24'b001111010100111101010111;
#1 $display("%b", po);
# 1  pi=24'b000100011010110010111001;
#1 $display("%b", po);
# 1  pi=24'b001010000101001100010111;
#1 $display("%b", po);
# 1  pi=24'b000010111100011000000011;
#1 $display("%b", po);
# 1  pi=24'b011001011011100110110101;
#1 $display("%b", po);
# 1  pi=24'b111110000100011011001010;
#1 $display("%b", po);
# 1  pi=24'b011100001101101100010001;
#1 $display("%b", po);
# 1  pi=24'b000101101001000000111111;
#1 $display("%b", po);
# 1  pi=24'b011101011011011101001010;
#1 $display("%b", po);
# 1  pi=24'b010111110110110100111011;
#1 $display("%b", po);
# 1  pi=24'b110100000101000110000001;
#1 $display("%b", po);
# 1  pi=24'b111011010000010010100111;
#1 $display("%b", po);
# 1  pi=24'b110101111000100110000101;
#1 $display("%b", po);
# 1  pi=24'b001110111010001101010110;
#1 $display("%b", po);
# 1  pi=24'b010000101100011000100011;
#1 $display("%b", po);
# 1  pi=24'b011110011111011011100010;
#1 $display("%b", po);
# 1  pi=24'b010010001100111100100111;
#1 $display("%b", po);
# 1  pi=24'b111110000101010101000100;
#1 $display("%b", po);
# 1  pi=24'b001110110111110010011011;
#1 $display("%b", po);
# 1  pi=24'b000000100110000100111010;
#1 $display("%b", po);
# 1  pi=24'b110001001000001010010100;
#1 $display("%b", po);
# 1  pi=24'b000010100011111010001000;
#1 $display("%b", po);
# 1  pi=24'b011100101001110000101110;
#1 $display("%b", po);
# 1  pi=24'b010110011000011111111010;
#1 $display("%b", po);
# 1  pi=24'b000001001011011100010110;
#1 $display("%b", po);
# 1  pi=24'b100011000101010110001010;
#1 $display("%b", po);
# 1  pi=24'b111010100010000000001101;
#1 $display("%b", po);
# 1  pi=24'b111110110110010001000110;
#1 $display("%b", po);
# 1  pi=24'b110010110000000111000111;
#1 $display("%b", po);
# 1  pi=24'b001001101000010111101000;
#1 $display("%b", po);
# 1  pi=24'b110011110011000110101001;
#1 $display("%b", po);
# 1  pi=24'b010001010110111110111111;
#1 $display("%b", po);
# 1  pi=24'b011011011110011111100110;
#1 $display("%b", po);
# 1  pi=24'b011110111100110010100101;
#1 $display("%b", po);
# 1  pi=24'b000111010110100001101010;
#1 $display("%b", po);
# 1  pi=24'b100111100001110101100011;
#1 $display("%b", po);
# 1  pi=24'b000000100000001110111101;
#1 $display("%b", po);
# 1  pi=24'b010011100100001111010011;
#1 $display("%b", po);
# 1  pi=24'b101111111110010111011101;
#1 $display("%b", po);
# 1  pi=24'b100101101101001000001110;
#1 $display("%b", po);
# 1  pi=24'b111111000110101000110011;
#1 $display("%b", po);
# 1  pi=24'b100101000110010111010101;
#1 $display("%b", po);
# 1  pi=24'b110001111101111011001111;
#1 $display("%b", po);
# 1  pi=24'b010000111110111000110111;
#1 $display("%b", po);
# 1  pi=24'b101000010010010110101001;
#1 $display("%b", po);
# 1  pi=24'b010100101000101011000001;
#1 $display("%b", po);
# 1  pi=24'b001111010101101110010010;
#1 $display("%b", po);
# 1  pi=24'b110011111110010001000101;
#1 $display("%b", po);
# 1  pi=24'b011100110101101111010001;
#1 $display("%b", po);
# 1  pi=24'b101010101011111101100011;
#1 $display("%b", po);
# 1  pi=24'b011010100011101100010110;
#1 $display("%b", po);
# 1  pi=24'b000010011110110110010111;
#1 $display("%b", po);
# 1  pi=24'b010001110001110110111010;
#1 $display("%b", po);
# 1  pi=24'b011111111011001001010000;
#1 $display("%b", po);
# 1  pi=24'b000011111111000110111100;
#1 $display("%b", po);
# 1  pi=24'b000100110000101000001010;
#1 $display("%b", po);
# 1  pi=24'b111101111000101000101110;
#1 $display("%b", po);
# 1  pi=24'b100000111010110011010111;
#1 $display("%b", po);
# 1  pi=24'b101100100100100110011100;
#1 $display("%b", po);
# 1  pi=24'b001110010101011010000001;
#1 $display("%b", po);
# 1  pi=24'b111111011110001111100000;
#1 $display("%b", po);
# 1  pi=24'b010000110011000101110100;
#1 $display("%b", po);
# 1  pi=24'b000010110101001100000110;
#1 $display("%b", po);
# 1  pi=24'b101110000001110001101011;
#1 $display("%b", po);
# 1  pi=24'b100011111011010100101110;
#1 $display("%b", po);
# 1  pi=24'b111001111010011000000010;
#1 $display("%b", po);
# 1  pi=24'b010011010011111110110010;
#1 $display("%b", po);
# 1  pi=24'b110110010011000011101001;
#1 $display("%b", po);
# 1  pi=24'b010110010100000011010010;
#1 $display("%b", po);
# 1  pi=24'b100100000110000110110110;
#1 $display("%b", po);
# 1  pi=24'b011100011111010100010011;
#1 $display("%b", po);
# 1  pi=24'b101011100011011111110011;
#1 $display("%b", po);
# 1  pi=24'b010010011101010001111101;
#1 $display("%b", po);
# 1  pi=24'b111010010100101110011111;
#1 $display("%b", po);
# 1  pi=24'b101100101011100010111101;
#1 $display("%b", po);
# 1  pi=24'b011011011000110000101010;
#1 $display("%b", po);
# 1  pi=24'b011101101111111010010001;
#1 $display("%b", po);
# 1  pi=24'b010110010101110110010001;
#1 $display("%b", po);
# 1  pi=24'b110011110110000010000001;
#1 $display("%b", po);
# 1  pi=24'b111011100010011000000110;
#1 $display("%b", po);
# 1  pi=24'b010010001011101000100111;
#1 $display("%b", po);
# 1  pi=24'b110001011000001111110110;
#1 $display("%b", po);
# 1  pi=24'b000011111011111100111110;
#1 $display("%b", po);
# 1  pi=24'b110000001001010001110110;
#1 $display("%b", po);
# 1  pi=24'b101111010111011110001001;
#1 $display("%b", po);
# 1  pi=24'b010010000101001101011110;
#1 $display("%b", po);
# 1  pi=24'b111011010100101011000101;
#1 $display("%b", po);
# 1  pi=24'b110000000010011011111110;
#1 $display("%b", po);
# 1  pi=24'b110110011010101011001000;
#1 $display("%b", po);
# 1  pi=24'b011101110110001001110001;
#1 $display("%b", po);
# 1  pi=24'b100111000011010100100101;
#1 $display("%b", po);
# 1  pi=24'b010000101101100001000011;
#1 $display("%b", po);
# 1  pi=24'b111100101011100100111011;
#1 $display("%b", po);
# 1  pi=24'b000010111000001101010011;
#1 $display("%b", po);
# 1  pi=24'b010011101000010001100110;
#1 $display("%b", po);
# 1  pi=24'b001001101010111000000110;
#1 $display("%b", po);
# 1  pi=24'b111000010000010101000110;
#1 $display("%b", po);
# 1  pi=24'b111111100101011011011011;
#1 $display("%b", po);
# 1  pi=24'b100010010100100011011011;
#1 $display("%b", po);
# 1  pi=24'b111101000010011111111000;
#1 $display("%b", po);
# 1  pi=24'b100010111111000110100011;
#1 $display("%b", po);
# 1  pi=24'b001100100001001111100100;
#1 $display("%b", po);
# 1  pi=24'b100110100011001100000100;
#1 $display("%b", po);
# 1  pi=24'b010100010000001111000100;
#1 $display("%b", po);
# 1  pi=24'b011001110100100110100011;
#1 $display("%b", po);
# 1  pi=24'b100010001011111001110111;
#1 $display("%b", po);
# 1  pi=24'b011101011011110100100000;
#1 $display("%b", po);
# 1  pi=24'b111000001101110100011001;
#1 $display("%b", po);
# 1  pi=24'b011000101100010101101111;
#1 $display("%b", po);
# 1  pi=24'b001010011110000010011110;
#1 $display("%b", po);
# 1  pi=24'b111101000001101101000100;
#1 $display("%b", po);
# 1  pi=24'b011101101111110101000111;
#1 $display("%b", po);
# 1  pi=24'b101001001000101100011101;
#1 $display("%b", po);
# 1  pi=24'b001000101001100110101001;
#1 $display("%b", po);
# 1  pi=24'b011111001000101000111001;
#1 $display("%b", po);
# 1  pi=24'b011101111000001100101000;
#1 $display("%b", po);
# 1  pi=24'b101100110000000001101001;
#1 $display("%b", po);
# 1  pi=24'b111111000011111101010011;
#1 $display("%b", po);
# 1  pi=24'b010011111001111011111011;
#1 $display("%b", po);
# 1  pi=24'b110001100010110001101111;
#1 $display("%b", po);
# 1  pi=24'b111100001000101010100110;
#1 $display("%b", po);
# 1  pi=24'b110000010101011101100011;
#1 $display("%b", po);
# 1  pi=24'b010110100010101011100100;
#1 $display("%b", po);
# 1  pi=24'b001100100110000101000110;
#1 $display("%b", po);
# 1  pi=24'b111101100111000001000000;
#1 $display("%b", po);
# 1  pi=24'b110111001011101011001001;
#1 $display("%b", po);
# 1  pi=24'b100001100111100111011100;
#1 $display("%b", po);
# 1  pi=24'b111001010110101101110110;
#1 $display("%b", po);
# 1  pi=24'b000010000011100100100001;
#1 $display("%b", po);
# 1  pi=24'b011010011100011101111101;
#1 $display("%b", po);
# 1  pi=24'b010000001111101110000111;
#1 $display("%b", po);
# 1  pi=24'b001111110010001011001001;
#1 $display("%b", po);
# 1  pi=24'b110000101111110110011010;
#1 $display("%b", po);
# 1  pi=24'b000001111101110110101011;
#1 $display("%b", po);
# 1  pi=24'b011100111101100101110000;
#1 $display("%b", po);
# 1  pi=24'b010110110001100001000010;
#1 $display("%b", po);
# 1  pi=24'b100000000001101011010101;
#1 $display("%b", po);
# 1  pi=24'b101000001100100010111111;
#1 $display("%b", po);
# 1  pi=24'b010100011000000011001011;
#1 $display("%b", po);
# 1  pi=24'b000100100011001111010101;
#1 $display("%b", po);
# 1  pi=24'b110100001001011101010100;
#1 $display("%b", po);
# 1  pi=24'b001000001010100001110011;
#1 $display("%b", po);
# 1  pi=24'b100010000111010111101100;
#1 $display("%b", po);
# 1  pi=24'b011111110010101000101010;
#1 $display("%b", po);
# 1  pi=24'b101010101101110011010001;
#1 $display("%b", po);
# 1  pi=24'b011101010110111001010010;
#1 $display("%b", po);
# 1  pi=24'b101101101000000101010111;
#1 $display("%b", po);
# 1  pi=24'b000001000100101001000001;
#1 $display("%b", po);
# 1  pi=24'b000000101010100001100001;
#1 $display("%b", po);
# 1  pi=24'b010011110010100010001101;
#1 $display("%b", po);
# 1  pi=24'b001000011110001010101101;
#1 $display("%b", po);
# 1  pi=24'b110111110000101110000001;
#1 $display("%b", po);
# 1  pi=24'b011001101001100111000011;
#1 $display("%b", po);
# 1  pi=24'b010110010000000011111100;
#1 $display("%b", po);
# 1  pi=24'b001001101100011011010011;
#1 $display("%b", po);
# 1  pi=24'b011000010011101000011000;
#1 $display("%b", po);
# 1  pi=24'b010000111101011001001000;
#1 $display("%b", po);
# 1  pi=24'b001101010011001110010010;
#1 $display("%b", po);
# 1  pi=24'b001100111001110010000111;
#1 $display("%b", po);
# 1  pi=24'b001011110001100111110110;
#1 $display("%b", po);
# 1  pi=24'b101110101100101101100001;
#1 $display("%b", po);
# 1  pi=24'b111110011100010000000011;
#1 $display("%b", po);
# 1  pi=24'b110111101010001011100000;
#1 $display("%b", po);
# 1  pi=24'b100100110011100111001101;
#1 $display("%b", po);
# 1  pi=24'b110100101011111010000110;
#1 $display("%b", po);
# 1  pi=24'b000001100000000001011000;
#1 $display("%b", po);
# 1  pi=24'b101010011001000110100010;
#1 $display("%b", po);
# 1  pi=24'b110000001101110000111010;
#1 $display("%b", po);
# 1  pi=24'b001011000101010010001110;
#1 $display("%b", po);
# 1  pi=24'b000110010111010001001011;
#1 $display("%b", po);
# 1  pi=24'b110011010100100111010011;
#1 $display("%b", po);
# 1  pi=24'b111101110000101000100001;
#1 $display("%b", po);
# 1  pi=24'b001000011000110100000000;
#1 $display("%b", po);
# 1  pi=24'b111111100111100110100100;
#1 $display("%b", po);
# 1  pi=24'b100110011001101110010101;
#1 $display("%b", po);
# 1  pi=24'b000111011001010001100011;
#1 $display("%b", po);
# 1  pi=24'b101011111100110011111000;
#1 $display("%b", po);
# 1  pi=24'b101011100001010110101111;
#1 $display("%b", po);
# 1  pi=24'b110101010010110101101001;
#1 $display("%b", po);
# 1  pi=24'b110010101000101000000000;
#1 $display("%b", po);
# 1  pi=24'b011001110100110111001101;
#1 $display("%b", po);
# 1  pi=24'b101011111010101111011010;
#1 $display("%b", po);
# 1  pi=24'b011110011001011001100010;
#1 $display("%b", po);
# 1  pi=24'b000001100011100001110100;
#1 $display("%b", po);
# 1  pi=24'b101000001011100101101110;
#1 $display("%b", po);
# 1  pi=24'b100110011110000111101011;
#1 $display("%b", po);
# 1  pi=24'b001001010101100010011110;
#1 $display("%b", po);
# 1  pi=24'b111010111111100110111001;
#1 $display("%b", po);
# 1  pi=24'b111110111010110101000010;
#1 $display("%b", po);
# 1  pi=24'b001110001011001110101111;
#1 $display("%b", po);
# 1  pi=24'b011100101101010100111011;
#1 $display("%b", po);
# 1  pi=24'b111100011010101101001010;
#1 $display("%b", po);
# 1  pi=24'b110000000100000110000010;
#1 $display("%b", po);
# 1  pi=24'b100111011001001010010100;
#1 $display("%b", po);
# 1  pi=24'b011110101010001101011111;
#1 $display("%b", po);
# 1  pi=24'b000111111011110011110001;
#1 $display("%b", po);
# 1  pi=24'b110110001000110101101101;
#1 $display("%b", po);
# 1  pi=24'b110110100001001101111001;
#1 $display("%b", po);
# 1  pi=24'b111111111000110111101010;
#1 $display("%b", po);
# 1  pi=24'b100111111111100110100011;
#1 $display("%b", po);
# 1  pi=24'b001100011110011001011001;
#1 $display("%b", po);
# 1  pi=24'b100001001001110000000101;
#1 $display("%b", po);
# 1  pi=24'b101011010011111000111010;
#1 $display("%b", po);
# 1  pi=24'b010001010010111111011001;
#1 $display("%b", po);
# 1  pi=24'b010100000001000111001110;
#1 $display("%b", po);
# 1  pi=24'b000000101111000100001001;
#1 $display("%b", po);
# 1  pi=24'b110011100101011111111101;
#1 $display("%b", po);
# 1  pi=24'b011101011001111100000011;
#1 $display("%b", po);
# 1  pi=24'b011010101110000101101111;
#1 $display("%b", po);
# 1  pi=24'b101111100101001110001101;
#1 $display("%b", po);
# 1  pi=24'b010100110011110000110100;
#1 $display("%b", po);
# 1  pi=24'b101010101000110001011001;
#1 $display("%b", po);
# 1  pi=24'b000010000111110110000000;
#1 $display("%b", po);
# 1  pi=24'b110110111010101101110100;
#1 $display("%b", po);
# 1  pi=24'b111110010011000000001100;
#1 $display("%b", po);
# 1  pi=24'b001110011000011110010110;
#1 $display("%b", po);
# 1  pi=24'b001110111000011000110001;
#1 $display("%b", po);
# 1  pi=24'b010101000101001010101111;
#1 $display("%b", po);
# 1  pi=24'b100011010100110001001111;
#1 $display("%b", po);
# 1  pi=24'b011000000100000001100011;
#1 $display("%b", po);
# 1  pi=24'b011111100110010011011011;
#1 $display("%b", po);
# 1  pi=24'b101010100011000101111100;
#1 $display("%b", po);
# 1  pi=24'b110010011100110100111100;
#1 $display("%b", po);
# 1  pi=24'b000010101010111001111111;
#1 $display("%b", po);
# 1  pi=24'b011010000111111010101010;
#1 $display("%b", po);
# 1  pi=24'b011001000000010001010100;
#1 $display("%b", po);
# 1  pi=24'b011000101101110010011110;
#1 $display("%b", po);
# 1  pi=24'b011011000000100001001101;
#1 $display("%b", po);
# 1  pi=24'b000010110111010011100000;
#1 $display("%b", po);
# 1  pi=24'b001111110111110100111111;
#1 $display("%b", po);
# 1  pi=24'b011001001010001111001110;
#1 $display("%b", po);
# 1  pi=24'b111000101100011010100011;
#1 $display("%b", po);
# 1  pi=24'b000001010110010100111001;
#1 $display("%b", po);
# 1  pi=24'b000010110001001110111010;
#1 $display("%b", po);
# 1  pi=24'b000100011111001000010001;
#1 $display("%b", po);
# 1  pi=24'b111100101101100001001110;
#1 $display("%b", po);
# 1  pi=24'b100000001110111110001101;
#1 $display("%b", po);
# 1  pi=24'b011001100100101000010001;
#1 $display("%b", po);
# 1  pi=24'b000110010011110111100111;
#1 $display("%b", po);
# 1  pi=24'b100000001110011101100111;
#1 $display("%b", po);
# 1  pi=24'b111010001110111100011001;
#1 $display("%b", po);
# 1  pi=24'b001100101010000011000100;
#1 $display("%b", po);
# 1  pi=24'b111101111100001101110001;
#1 $display("%b", po);
# 1  pi=24'b111111000111100010111110;
#1 $display("%b", po);
# 1  pi=24'b011000011110101101111110;
#1 $display("%b", po);
# 1  pi=24'b001101011001101010011010;
#1 $display("%b", po);
# 1  pi=24'b011011001000001110101111;
#1 $display("%b", po);
# 1  pi=24'b100111011110011000011010;
#1 $display("%b", po);
# 1  pi=24'b100111100111100100110011;
#1 $display("%b", po);
# 1  pi=24'b010000001111000010100001;
#1 $display("%b", po);
# 1  pi=24'b100100111010011100000011;
#1 $display("%b", po);
# 1  pi=24'b100111011101001100100110;
#1 $display("%b", po);
# 1  pi=24'b001011110010000101111100;
#1 $display("%b", po);
# 1  pi=24'b000000100101110010100000;
#1 $display("%b", po);
# 1  pi=24'b010011110001011000100110;
#1 $display("%b", po);
# 1  pi=24'b111011110011110110100011;
#1 $display("%b", po);
# 1  pi=24'b001110000111101111001100;
#1 $display("%b", po);
# 1  pi=24'b010011001101000000111111;
#1 $display("%b", po);
# 1  pi=24'b010010110001001110111101;
#1 $display("%b", po);
# 1  pi=24'b010101010000111001010011;
#1 $display("%b", po);
# 1  pi=24'b100100010010110001010010;
#1 $display("%b", po);
# 1  pi=24'b010101110010101011011001;
#1 $display("%b", po);
# 1  pi=24'b001001010011001100100000;
#1 $display("%b", po);
# 1  pi=24'b000010111010000100110001;
#1 $display("%b", po);
# 1  pi=24'b100010011100100001110011;
#1 $display("%b", po);
# 1  pi=24'b000110100100001101111101;
#1 $display("%b", po);
# 1  pi=24'b101111111001110000010111;
#1 $display("%b", po);
# 1  pi=24'b101101010111011011001001;
#1 $display("%b", po);
# 1  pi=24'b010111000110111110001101;
#1 $display("%b", po);
# 1  pi=24'b010110010101010011110100;
#1 $display("%b", po);
# 1  pi=24'b110101110010100011010100;
#1 $display("%b", po);
# 1  pi=24'b101110010000111101101101;
#1 $display("%b", po);
# 1  pi=24'b110011010110001011000101;
#1 $display("%b", po);
# 1  pi=24'b110000111101111010001000;
#1 $display("%b", po);
# 1  pi=24'b100100010110011100010011;
#1 $display("%b", po);
# 1  pi=24'b100100100001100111100010;
#1 $display("%b", po);
# 1  pi=24'b111001110011100001010111;
#1 $display("%b", po);
# 1  pi=24'b011111111011001110110100;
#1 $display("%b", po);
# 1  pi=24'b100001101000101100101011;
#1 $display("%b", po);
# 1  pi=24'b000111101101110111001111;
#1 $display("%b", po);
# 1  pi=24'b011011100010000001011100;
#1 $display("%b", po);
# 1  pi=24'b001111001001000001011000;
#1 $display("%b", po);
# 1  pi=24'b101110011110000010110011;
#1 $display("%b", po);
# 1  pi=24'b001001001100001111100111;
#1 $display("%b", po);
# 1  pi=24'b010000111000011011100001;
#1 $display("%b", po);
# 1  pi=24'b010111111011000000110110;
#1 $display("%b", po);
# 1  pi=24'b111101000000001111100100;
#1 $display("%b", po);
# 1  pi=24'b101110001110101011000001;
#1 $display("%b", po);
# 1  pi=24'b001010000010000110101110;
#1 $display("%b", po);
# 1  pi=24'b011101101101111111011100;
#1 $display("%b", po);
# 1  pi=24'b100010000011000100000000;
#1 $display("%b", po);
# 1  pi=24'b010111100000011000001011;
#1 $display("%b", po);
# 1  pi=24'b100001001101011001101100;
#1 $display("%b", po);
# 1  pi=24'b011000010011101101110110;
#1 $display("%b", po);
# 1  pi=24'b000110100110010010101000;
#1 $display("%b", po);
# 1  pi=24'b001001100010100000101100;
#1 $display("%b", po);
# 1  pi=24'b000011011101101110111110;
#1 $display("%b", po);
# 1  pi=24'b010000111111110001101010;
#1 $display("%b", po);
# 1  pi=24'b010011001100101011001001;
#1 $display("%b", po);
# 1  pi=24'b101000010001000010110111;
#1 $display("%b", po);
# 1  pi=24'b110010010110111011011001;
#1 $display("%b", po);
# 1  pi=24'b000011000011011110001010;
#1 $display("%b", po);
# 1  pi=24'b000101010011111010100100;
#1 $display("%b", po);
# 1  pi=24'b111110110010111111100110;
#1 $display("%b", po);
# 1  pi=24'b010111111110110101111001;
#1 $display("%b", po);
# 1  pi=24'b001000010110101011101101;
#1 $display("%b", po);
# 1  pi=24'b011110000000110111000100;
#1 $display("%b", po);
# 1  pi=24'b011110001011110101110100;
#1 $display("%b", po);
# 1  pi=24'b111010000000011000001111;
#1 $display("%b", po);
# 1  pi=24'b111111011000110000110011;
#1 $display("%b", po);
# 1  pi=24'b011011001011110110100010;
#1 $display("%b", po);
# 1  pi=24'b110110101100110111010111;
#1 $display("%b", po);
# 1  pi=24'b101010000000000111010100;
#1 $display("%b", po);
# 1  pi=24'b111011110101110101111010;
#1 $display("%b", po);
# 1  pi=24'b110101101001001101001100;
#1 $display("%b", po);
# 1  pi=24'b011001011111110010010110;
#1 $display("%b", po);
# 1  pi=24'b100101010010011111110110;
#1 $display("%b", po);
# 1  pi=24'b010100010110000101100001;
#1 $display("%b", po);
# 1  pi=24'b111101100001000111001000;
#1 $display("%b", po);
# 1  pi=24'b110001001001001010101101;
#1 $display("%b", po);
# 1  pi=24'b101000010110001111001011;
#1 $display("%b", po);
# 1  pi=24'b010000100000000110110011;
#1 $display("%b", po);
# 1  pi=24'b000100010110000001010001;
#1 $display("%b", po);
# 1  pi=24'b010111101011100110111101;
#1 $display("%b", po);
# 1  pi=24'b000011010100010110000011;
#1 $display("%b", po);
# 1  pi=24'b100011011000100101000101;
#1 $display("%b", po);
# 1  pi=24'b001110010011010001010010;
#1 $display("%b", po);
# 1  pi=24'b001110010000111001001100;
#1 $display("%b", po);
# 1  pi=24'b100000110101111111101100;
#1 $display("%b", po);
# 1  pi=24'b011100101010100111010101;
#1 $display("%b", po);
# 1  pi=24'b100111010010001000110111;
#1 $display("%b", po);
# 1  pi=24'b111000111111000000000101;
#1 $display("%b", po);
# 1  pi=24'b000111001101100001010000;
#1 $display("%b", po);
# 1  pi=24'b110101111101100101110100;
#1 $display("%b", po);
# 1  pi=24'b000001011110101000001110;
#1 $display("%b", po);
# 1  pi=24'b111101101010010111101101;
#1 $display("%b", po);
# 1  pi=24'b110111111000010110110101;
#1 $display("%b", po);
# 1  pi=24'b000101110011100101100011;
#1 $display("%b", po);
# 1  pi=24'b110000001100000001011011;
#1 $display("%b", po);
# 1  pi=24'b000111101001101001010111;
#1 $display("%b", po);
# 1  pi=24'b001101010010010101011101;
#1 $display("%b", po);
# 1  pi=24'b001111111100010000010000;
#1 $display("%b", po);
# 1  pi=24'b101101101100010100001101;
#1 $display("%b", po);
# 1  pi=24'b111011101001010100111010;
#1 $display("%b", po);
# 1  pi=24'b010000010010110010001111;
#1 $display("%b", po);
# 1  pi=24'b001110101010011101111100;
#1 $display("%b", po);
# 1  pi=24'b101010011110000011011010;
#1 $display("%b", po);
# 1  pi=24'b111111110000110111111101;
#1 $display("%b", po);
# 1  pi=24'b000101100111011110111111;
#1 $display("%b", po);
# 1  pi=24'b111110011001110100110111;
#1 $display("%b", po);
# 1  pi=24'b010111001000010010000100;
#1 $display("%b", po);
# 1  pi=24'b000101101011001010110100;
#1 $display("%b", po);
# 1  pi=24'b101101111000000110101100;
#1 $display("%b", po);
# 1  pi=24'b100100010101001101000010;
#1 $display("%b", po);
# 1  pi=24'b100011111010100001100010;
#1 $display("%b", po);
# 1  pi=24'b011011101001001100000100;
#1 $display("%b", po);
# 1  pi=24'b000011111110100100000010;
#1 $display("%b", po);
# 1  pi=24'b101001010011011010010001;
#1 $display("%b", po);
# 1  pi=24'b001011101101111100101001;
#1 $display("%b", po);
# 1  pi=24'b010100101100011010101000;
#1 $display("%b", po);
# 1  pi=24'b111111101101001001010000;
#1 $display("%b", po);
# 1  pi=24'b000101010010110100000100;
#1 $display("%b", po);
# 1  pi=24'b111100010111010001010000;
#1 $display("%b", po);
# 1  pi=24'b000101011111010010110001;
#1 $display("%b", po);
# 1  pi=24'b010111110101010011110100;
#1 $display("%b", po);
# 1  pi=24'b011110111001000100010110;
#1 $display("%b", po);
# 1  pi=24'b000000100001011111010100;
#1 $display("%b", po);
# 1  pi=24'b001010110011100100011011;
#1 $display("%b", po);
# 1  pi=24'b101001110000010100101100;
#1 $display("%b", po);
# 1  pi=24'b101101000000111001100111;
#1 $display("%b", po);
# 1  pi=24'b010001111001111010000000;
#1 $display("%b", po);
# 1  pi=24'b100101001100111011100010;
#1 $display("%b", po);
# 1  pi=24'b100000110001110011001101;
#1 $display("%b", po);
# 1  pi=24'b101110001010111101000011;
#1 $display("%b", po);
# 1  pi=24'b001000010000011111100000;
#1 $display("%b", po);
# 1  pi=24'b000101000101001000001011;
#1 $display("%b", po);
# 1  pi=24'b101110000111110111000110;
#1 $display("%b", po);
# 1  pi=24'b000110110110010110001011;
#1 $display("%b", po);
# 1  pi=24'b000000001011010100110001;
#1 $display("%b", po);
# 1  pi=24'b110000000110101101111011;
#1 $display("%b", po);
# 1  pi=24'b001000001101010101010011;
#1 $display("%b", po);
# 1  pi=24'b000110111100000000010100;
#1 $display("%b", po);
# 1  pi=24'b110101111010100001101101;
#1 $display("%b", po);
# 1  pi=24'b000011001000100000111101;
#1 $display("%b", po);
# 1  pi=24'b000010001000010010000011;
#1 $display("%b", po);
# 1  pi=24'b101000101100111011100101;
#1 $display("%b", po);
# 1  pi=24'b111110101000000000010011;
#1 $display("%b", po);
# 1  pi=24'b001000100010101000000111;
#1 $display("%b", po);
# 1  pi=24'b111111000101010111011110;
#1 $display("%b", po);
# 1  pi=24'b001100000111011101001011;
#1 $display("%b", po);
# 1  pi=24'b110100011010001110000101;
#1 $display("%b", po);
# 1  pi=24'b100000000010010111000011;
#1 $display("%b", po);
# 1  pi=24'b010111001010101101000110;
#1 $display("%b", po);
# 1  pi=24'b101101011010011000110101;
#1 $display("%b", po);
# 1  pi=24'b000000011101000010110010;
#1 $display("%b", po);
# 1  pi=24'b111010100000100010011000;
#1 $display("%b", po);
# 1  pi=24'b111010100101100110011010;
#1 $display("%b", po);
# 1  pi=24'b011100110101000011110110;
#1 $display("%b", po);
# 1  pi=24'b001001000001000001101000;
#1 $display("%b", po);
# 1  pi=24'b111011100101000111101000;
#1 $display("%b", po);
# 1  pi=24'b100000001011000001101100;
#1 $display("%b", po);
# 1  pi=24'b111001000111100110011010;
#1 $display("%b", po);
# 1  pi=24'b111111111001110001111101;
#1 $display("%b", po);
# 1  pi=24'b110001101110001001000010;
#1 $display("%b", po);
# 1  pi=24'b110111010001101000011010;
#1 $display("%b", po);
# 1  pi=24'b010100011110110000011101;
#1 $display("%b", po);
# 1  pi=24'b100101011101100011000000;
#1 $display("%b", po);
# 1  pi=24'b101000100010100000011010;
#1 $display("%b", po);
# 1  pi=24'b001101001110100001111100;
#1 $display("%b", po);
# 1  pi=24'b011011010111111100001110;
#1 $display("%b", po);
# 1  pi=24'b001101011010011000100111;
#1 $display("%b", po);
# 1  pi=24'b011010101010000110100100;
#1 $display("%b", po);
# 1  pi=24'b101111000100011011000111;
#1 $display("%b", po);
# 1  pi=24'b010100000111000110011010;
#1 $display("%b", po);
# 1  pi=24'b100010000111000010011011;
#1 $display("%b", po);
# 1  pi=24'b011101111101101101000010;
#1 $display("%b", po);
# 1  pi=24'b111110011000100110000110;
#1 $display("%b", po);
# 1  pi=24'b000010110010111000101010;
#1 $display("%b", po);
# 1  pi=24'b011001000001110011100111;
#1 $display("%b", po);
# 1  pi=24'b001001010010100000110110;
#1 $display("%b", po);
# 1  pi=24'b001001101110010011001110;
#1 $display("%b", po);
# 1  pi=24'b000101110010001011001000;
#1 $display("%b", po);
# 1  pi=24'b000010010110110000100111;
#1 $display("%b", po);
# 1  pi=24'b101000000011010010001111;
#1 $display("%b", po);
# 1  pi=24'b010010000000011000100111;
#1 $display("%b", po);
# 1  pi=24'b111000111011000111001001;
#1 $display("%b", po);
# 1  pi=24'b111010111011111101110101;
#1 $display("%b", po);
# 1  pi=24'b011000111000110010010011;
#1 $display("%b", po);
# 1  pi=24'b100000110010000001100110;
#1 $display("%b", po);
# 1  pi=24'b110010001010110110011111;
#1 $display("%b", po);
# 1  pi=24'b001000011010010111100111;
#1 $display("%b", po);
# 1  pi=24'b011110101011100000011100;
#1 $display("%b", po);
# 1  pi=24'b011001111100001000101010;
#1 $display("%b", po);
# 1  pi=24'b001111100000010010110011;
#1 $display("%b", po);
# 1  pi=24'b000110011011111010010011;
#1 $display("%b", po);
# 1  pi=24'b000000010110100111100010;
#1 $display("%b", po);
# 1  pi=24'b010100100011100111100111;
#1 $display("%b", po);
# 1  pi=24'b110011000000111100010111;
#1 $display("%b", po);
# 1  pi=24'b101000001001000100001100;
#1 $display("%b", po);
# 1  pi=24'b100010100001110101010100;
#1 $display("%b", po);
# 1  pi=24'b010110110100100001011000;
#1 $display("%b", po);
# 1  pi=24'b000001101001010110110011;
#1 $display("%b", po);
# 1  pi=24'b010110101001100011100001;
#1 $display("%b", po);
# 1  pi=24'b011101101101101010010100;
#1 $display("%b", po);
# 1  pi=24'b100001000011000111011100;
#1 $display("%b", po);
# 1  pi=24'b001100001000100101100001;
#1 $display("%b", po);
# 1  pi=24'b001000001100001001000001;
#1 $display("%b", po);
# 1  pi=24'b100001101010011000010000;
#1 $display("%b", po);
# 1  pi=24'b101011011100001101011100;
#1 $display("%b", po);
# 1  pi=24'b010100010101010110111011;
#1 $display("%b", po);
# 1  pi=24'b111110010011101100011101;
#1 $display("%b", po);
# 1  pi=24'b110100010010010111011000;
#1 $display("%b", po);
# 1  pi=24'b001001110111100110001001;
#1 $display("%b", po);
# 1  pi=24'b010100110001000101010111;
#1 $display("%b", po);
# 1  pi=24'b010100001110110100101010;
#1 $display("%b", po);
# 1  pi=24'b001110011101111011111111;
#1 $display("%b", po);
# 1  pi=24'b010010100100111010100010;
#1 $display("%b", po);
# 1  pi=24'b011010101000010000100000;
#1 $display("%b", po);
# 1  pi=24'b110000001001011000001101;
#1 $display("%b", po);
# 1  pi=24'b011100100000111010001001;
#1 $display("%b", po);
# 1  pi=24'b000110000101110100100001;
#1 $display("%b", po);
# 1  pi=24'b100100101000110111001010;
#1 $display("%b", po);
# 1  pi=24'b111010100010111110100011;
#1 $display("%b", po);
# 1  pi=24'b010001100000000011110100;
#1 $display("%b", po);
# 1  pi=24'b101111110000011110110011;
#1 $display("%b", po);
# 1  pi=24'b011110000000101110010111;
#1 $display("%b", po);
# 1  pi=24'b011010011011110111101000;
#1 $display("%b", po);
# 1  pi=24'b100110001100110011111000;
#1 $display("%b", po);
# 1  pi=24'b111100111011000101011011;
#1 $display("%b", po);
# 1  pi=24'b111001110011000000110000;
#1 $display("%b", po);
# 1  pi=24'b001111101100011000010000;
#1 $display("%b", po);
# 1  pi=24'b110111000000000010110100;
#1 $display("%b", po);
# 1  pi=24'b101100110000011000001000;
#1 $display("%b", po);
# 1  pi=24'b101101001011000110010110;
#1 $display("%b", po);
# 1  pi=24'b110000011010111010000001;
#1 $display("%b", po);
# 1  pi=24'b011001101110111101010110;
#1 $display("%b", po);
# 1  pi=24'b101110010010010111110101;
#1 $display("%b", po);
# 1  pi=24'b001101000010111001100010;
#1 $display("%b", po);
# 1  pi=24'b001011111010110011100111;
#1 $display("%b", po);
# 1  pi=24'b000101001011110011011011;
#1 $display("%b", po);
# 1  pi=24'b011101100100010111100010;
#1 $display("%b", po);
# 1  pi=24'b001010111001011110101001;
#1 $display("%b", po);
# 1  pi=24'b010011110011000000100011;
#1 $display("%b", po);
# 1  pi=24'b110110101010000100001011;
#1 $display("%b", po);
# 1  pi=24'b101100001001010100000001;
#1 $display("%b", po);
# 1  pi=24'b101000011001111101001010;
#1 $display("%b", po);
# 1  pi=24'b011000100111110011010101;
#1 $display("%b", po);
# 1  pi=24'b111100101111010010100111;
#1 $display("%b", po);
# 1  pi=24'b110001101010101001001001;
#1 $display("%b", po);
# 1  pi=24'b101100001110011001001010;
#1 $display("%b", po);
# 1  pi=24'b000001001011011101010100;
#1 $display("%b", po);
# 1  pi=24'b101010101010000101110011;
#1 $display("%b", po);
# 1  pi=24'b010101111000011010101111;
#1 $display("%b", po);
# 1  pi=24'b001010011100000110010001;
#1 $display("%b", po);
# 1  pi=24'b000100111001100001001111;
#1 $display("%b", po);
# 1  pi=24'b100100101101111101100011;
#1 $display("%b", po);
# 1  pi=24'b100111010000010010010111;
#1 $display("%b", po);
# 1  pi=24'b010110100101111001100111;
#1 $display("%b", po);
# 1  pi=24'b010111000101110011011001;
#1 $display("%b", po);
# 1  pi=24'b001011010111010001100100;
#1 $display("%b", po);
# 1  pi=24'b011110110000111001101000;
#1 $display("%b", po);
# 1  pi=24'b001100000111011110100011;
#1 $display("%b", po);
# 1  pi=24'b001011010111101001101001;
#1 $display("%b", po);
# 1  pi=24'b001000011100101101100100;
#1 $display("%b", po);
# 1  pi=24'b000110111100001101110110;
#1 $display("%b", po);
# 1  pi=24'b101111011111001111000111;
#1 $display("%b", po);
# 1  pi=24'b000000010000001111001111;
#1 $display("%b", po);
# 1  pi=24'b000001010001011111110000;
#1 $display("%b", po);
# 1  pi=24'b001010001011111000111110;
#1 $display("%b", po);
# 1  pi=24'b010011000101100100011110;
#1 $display("%b", po);
# 1  pi=24'b110101101101100101000001;
#1 $display("%b", po);
# 1  pi=24'b111001100001001011110101;
#1 $display("%b", po);
# 1  pi=24'b010110001100010100001001;
#1 $display("%b", po);
# 1  pi=24'b100011011001011010010101;
#1 $display("%b", po);
# 1  pi=24'b101101000111010111010000;
#1 $display("%b", po);
# 1  pi=24'b100111111100001001111010;
#1 $display("%b", po);
# 1  pi=24'b010001111010001101111110;
#1 $display("%b", po);
# 1  pi=24'b000010001000011010000000;
#1 $display("%b", po);
# 1  pi=24'b011010001110101101011000;
#1 $display("%b", po);
# 1  pi=24'b010011011110100110111100;
#1 $display("%b", po);
# 1  pi=24'b000111010000101001001111;
#1 $display("%b", po);
# 1  pi=24'b111000111110100010111000;
#1 $display("%b", po);
# 1  pi=24'b000001111011100110011011;
#1 $display("%b", po);
# 1  pi=24'b111101001101111010111001;
#1 $display("%b", po);
# 1  pi=24'b011001101001000100101011;
#1 $display("%b", po);
# 1  pi=24'b111111101111110110011100;
#1 $display("%b", po);
# 1  pi=24'b111100001110100110000000;
#1 $display("%b", po);
# 1  pi=24'b010001011011010101000100;
#1 $display("%b", po);
# 1  pi=24'b001000010100010111100010;
#1 $display("%b", po);
# 1  pi=24'b011101111111011001100010;
#1 $display("%b", po);
# 1  pi=24'b111110010000011111000101;
#1 $display("%b", po);
# 1  pi=24'b110110111101010010000110;
#1 $display("%b", po);
# 1  pi=24'b111100100110100100101011;
#1 $display("%b", po);
# 1  pi=24'b001011111011110111100111;
#1 $display("%b", po);
# 1  pi=24'b010111111010011101001110;
#1 $display("%b", po);
# 1  pi=24'b110011000000011000001111;
#1 $display("%b", po);
# 1  pi=24'b011001010010110101000110;
#1 $display("%b", po);
# 1  pi=24'b011111000000001011001010;
#1 $display("%b", po);
# 1  pi=24'b111011100001011111110101;
#1 $display("%b", po);
# 1  pi=24'b001000010111100110110111;
#1 $display("%b", po);
# 1  pi=24'b001101110110000111101100;
#1 $display("%b", po);
# 1  pi=24'b011000111000011101101110;
#1 $display("%b", po);
# 1  pi=24'b111011110000000011010101;
#1 $display("%b", po);
# 1  pi=24'b000010101111000111001100;
#1 $display("%b", po);
# 1  pi=24'b100000100010001101001001;
#1 $display("%b", po);
# 1  pi=24'b001101010001001000111010;
#1 $display("%b", po);
# 1  pi=24'b111100011111010010100011;
#1 $display("%b", po);
# 1  pi=24'b110000000011110011000011;
#1 $display("%b", po);
# 1  pi=24'b101100001110111100111011;
#1 $display("%b", po);
# 1  pi=24'b011110100000001011010001;
#1 $display("%b", po);
# 1  pi=24'b101100101000000110110010;
#1 $display("%b", po);
# 1  pi=24'b110011101110001110110000;
#1 $display("%b", po);
# 1  pi=24'b100110100001111110101011;
#1 $display("%b", po);
# 1  pi=24'b100111000010110000001001;
#1 $display("%b", po);
# 1  pi=24'b000010011100101100011010;
#1 $display("%b", po);
# 1  pi=24'b000110000010100010101110;
#1 $display("%b", po);
# 1  pi=24'b100110000000111101101010;
#1 $display("%b", po);
# 1  pi=24'b011001000010011011010100;
#1 $display("%b", po);
# 1  pi=24'b000000010011111000010011;
#1 $display("%b", po);
# 1  pi=24'b010110100011010010101100;
#1 $display("%b", po);
# 1  pi=24'b100100111001000010111000;
#1 $display("%b", po);
# 1  pi=24'b001011110001010101001100;
#1 $display("%b", po);
# 1  pi=24'b110000110001011101111001;
#1 $display("%b", po);
# 1  pi=24'b110011111110001111101101;
#1 $display("%b", po);
# 1  pi=24'b100000100101110111000111;
#1 $display("%b", po);
# 1  pi=24'b010111110111011100011100;
#1 $display("%b", po);
# 1  pi=24'b100000111001101111000101;
#1 $display("%b", po);
# 1  pi=24'b111110101101100100000001;
#1 $display("%b", po);
# 1  pi=24'b111001101001101001011000;
#1 $display("%b", po);
# 1  pi=24'b011110100101110100100110;
#1 $display("%b", po);
# 1  pi=24'b110000001101000000110001;
#1 $display("%b", po);
# 1  pi=24'b000111111101111000110001;
#1 $display("%b", po);
# 1  pi=24'b111111000011010111001110;
#1 $display("%b", po);
# 1  pi=24'b000101111001011000110010;
#1 $display("%b", po);
# 1  pi=24'b011000110011111110100111;
#1 $display("%b", po);
# 1  pi=24'b000100110111000000111001;
#1 $display("%b", po);
# 1  pi=24'b010000011011111010010001;
#1 $display("%b", po);
# 1  pi=24'b011010110000110011001011;
#1 $display("%b", po);
# 1  pi=24'b110010101101100100101110;
#1 $display("%b", po);
# 1  pi=24'b100001100101101010100100;
#1 $display("%b", po);
# 1  pi=24'b101011010010111101000000;
#1 $display("%b", po);
# 1  pi=24'b000010111101111110110001;
#1 $display("%b", po);
# 1  pi=24'b001000101011110110000100;
#1 $display("%b", po);
# 1  pi=24'b011001100101010110000101;
#1 $display("%b", po);
# 1  pi=24'b010011101100111001101011;
#1 $display("%b", po);
# 1  pi=24'b011000110011000000000011;
#1 $display("%b", po);
# 1  pi=24'b000110110001110011001111;
#1 $display("%b", po);
# 1  pi=24'b010101001111100110011101;
#1 $display("%b", po);
# 1  pi=24'b001011101101001101000110;
#1 $display("%b", po);
# 1  pi=24'b111101011111010011110001;
#1 $display("%b", po);
# 1  pi=24'b010101100111011000001101;
#1 $display("%b", po);
# 1  pi=24'b110111001010100110100000;
#1 $display("%b", po);
# 1  pi=24'b011010111001001011110001;
#1 $display("%b", po);
# 1  pi=24'b110110111101110011010110;
#1 $display("%b", po);
# 1  pi=24'b101011100001001100011011;
#1 $display("%b", po);
# 1  pi=24'b101100101000000100110110;
#1 $display("%b", po);
# 1  pi=24'b110110101111110011110000;
#1 $display("%b", po);
# 1  pi=24'b101110011111010101101110;
#1 $display("%b", po);
# 1  pi=24'b010110000001010000001010;
#1 $display("%b", po);
# 1  pi=24'b100001001010000011110001;
#1 $display("%b", po);
# 1  pi=24'b001111011010101000111100;
#1 $display("%b", po);
# 1  pi=24'b110011001010100111001111;
#1 $display("%b", po);
# 1  pi=24'b010001010010111011000010;
#1 $display("%b", po);
# 1  pi=24'b110000000111011101010110;
#1 $display("%b", po);
# 1  pi=24'b010001000011110110001010;
#1 $display("%b", po);
# 1  pi=24'b110000000011101010001110;
#1 $display("%b", po);
# 1  pi=24'b111000110001101001111101;
#1 $display("%b", po);
# 1  pi=24'b011000011010100110101111;
#1 $display("%b", po);
# 1  pi=24'b011100000010010111011100;
#1 $display("%b", po);
# 1  pi=24'b110010000100100001101010;
#1 $display("%b", po);
# 1  pi=24'b111001101101111000001110;
#1 $display("%b", po);
# 1  pi=24'b100001110010100011001100;
#1 $display("%b", po);
# 1  pi=24'b000100100000101000111000;
#1 $display("%b", po);
# 1  pi=24'b111001111110101110111011;
#1 $display("%b", po);
# 1  pi=24'b111101111011101011110111;
#1 $display("%b", po);
# 1  pi=24'b001010011000010100010001;
#1 $display("%b", po);
# 1  pi=24'b011001011100011011011001;
#1 $display("%b", po);
# 1  pi=24'b000000010110111110011001;
#1 $display("%b", po);
# 1  pi=24'b001111001101001100010111;
#1 $display("%b", po);
# 1  pi=24'b011100101100011101101110;
#1 $display("%b", po);
# 1  pi=24'b110111111101011000111101;
#1 $display("%b", po);
# 1  pi=24'b110000101010101111011100;
#1 $display("%b", po);
# 1  pi=24'b011001101001001111000001;
#1 $display("%b", po);
# 1  pi=24'b000010001000110001000111;
#1 $display("%b", po);
# 1  pi=24'b001111100010010101011110;
#1 $display("%b", po);
# 1  pi=24'b011101111001101101100010;
#1 $display("%b", po);
# 1  pi=24'b010111100010001101011100;
#1 $display("%b", po);
# 1  pi=24'b011101001001111000101001;
#1 $display("%b", po);
# 1  pi=24'b001110100111110100100011;
#1 $display("%b", po);
# 1  pi=24'b101100100011010011010111;
#1 $display("%b", po);
# 1  pi=24'b100011011010000001101111;
#1 $display("%b", po);
# 1  pi=24'b000011110001010110100011;
#1 $display("%b", po);
# 1  pi=24'b010010111001100110110111;
#1 $display("%b", po);
# 1  pi=24'b100001010110010100100100;
#1 $display("%b", po);
# 1  pi=24'b011101000111010101000100;
#1 $display("%b", po);
# 1  pi=24'b110001000001100001010100;
#1 $display("%b", po);
# 1  pi=24'b000110000100000101110001;
#1 $display("%b", po);
# 1  pi=24'b100000111100010001101111;
#1 $display("%b", po);
# 1  pi=24'b110101001001111111001000;
#1 $display("%b", po);
# 1  pi=24'b001101101111001010111100;
#1 $display("%b", po);
# 1  pi=24'b111101001000001101100100;
#1 $display("%b", po);
# 1  pi=24'b011101111101011101010100;
#1 $display("%b", po);
# 1  pi=24'b100000100001111110110010;
#1 $display("%b", po);
# 1  pi=24'b010101100001100001000010;
#1 $display("%b", po);
# 1  pi=24'b111001111010001111110110;
#1 $display("%b", po);
# 1  pi=24'b000010011011001111100010;
#1 $display("%b", po);
# 1  pi=24'b110110100100000000000110;
#1 $display("%b", po);
# 1  pi=24'b000100000011111011111101;
#1 $display("%b", po);
# 1  pi=24'b111000000010010000011001;
#1 $display("%b", po);
# 1  pi=24'b111000010000100000000001;
#1 $display("%b", po);
# 1  pi=24'b111100110010100011001100;
#1 $display("%b", po);
# 1  pi=24'b101101000101010011101011;
#1 $display("%b", po);
# 1  pi=24'b000010010011000010011110;
#1 $display("%b", po);
# 1  pi=24'b000010011010101110000100;
#1 $display("%b", po);
# 1  pi=24'b010111011100000100110100;
#1 $display("%b", po);
# 1  pi=24'b010010010101100101001000;
#1 $display("%b", po);
# 1  pi=24'b111011011101001011000001;
#1 $display("%b", po);
# 1  pi=24'b000110011011011010101001;
#1 $display("%b", po);
# 1  pi=24'b110001000000101110100000;
#1 $display("%b", po);
# 1  pi=24'b001111101101111000111000;
#1 $display("%b", po);
# 1  pi=24'b011110010110101101000110;
#1 $display("%b", po);
# 1  pi=24'b010010000100101111001101;
#1 $display("%b", po);
# 1  pi=24'b000100000011001100000100;
#1 $display("%b", po);
# 1  pi=24'b011000101101000001100101;
#1 $display("%b", po);
# 1  pi=24'b111110100001000111000011;
#1 $display("%b", po);
# 1  pi=24'b111100111011111101111100;
#1 $display("%b", po);
# 1  pi=24'b101101110001011101110110;
#1 $display("%b", po);
# 1  pi=24'b111011101000101010011001;
#1 $display("%b", po);
# 1  pi=24'b010010011001001110100011;
#1 $display("%b", po);
# 1  pi=24'b111011001010010011001101;
#1 $display("%b", po);
# 1  pi=24'b101010101100001111001010;
#1 $display("%b", po);
# 1  pi=24'b111111010001001100001100;
#1 $display("%b", po);
# 1  pi=24'b010000100101001101101010;
#1 $display("%b", po);
# 1  pi=24'b001000011110011111011100;
#1 $display("%b", po);
# 1  pi=24'b001110010011101110010010;
#1 $display("%b", po);
# 1  pi=24'b100101011001011000001101;
#1 $display("%b", po);
# 1  pi=24'b001110001000011010001100;
#1 $display("%b", po);
# 1  pi=24'b011100111000000011010001;
#1 $display("%b", po);
# 1  pi=24'b111010000101111011010000;
#1 $display("%b", po);
# 1  pi=24'b011010010100110110011101;
#1 $display("%b", po);
# 1  pi=24'b111110111000010101010011;
#1 $display("%b", po);
# 1  pi=24'b110110110111110000110000;
#1 $display("%b", po);
# 1  pi=24'b000001110011100100000110;
#1 $display("%b", po);
# 1  pi=24'b000001001100011000100001;
#1 $display("%b", po);
# 1  pi=24'b101011101100110010100001;
#1 $display("%b", po);
# 1  pi=24'b000001010001101010011100;
#1 $display("%b", po);
# 1  pi=24'b110001111000001011111110;
#1 $display("%b", po);
# 1  pi=24'b110010010101100100100111;
#1 $display("%b", po);
# 1  pi=24'b000100000001101110000100;
#1 $display("%b", po);
# 1  pi=24'b100111110100111100001010;
#1 $display("%b", po);
# 1  pi=24'b111010110011101111101001;
#1 $display("%b", po);
# 1  pi=24'b101001101011110111001010;
#1 $display("%b", po);
# 1  pi=24'b110000111011110001011001;
#1 $display("%b", po);
# 1  pi=24'b001101110101110001010000;
#1 $display("%b", po);
# 1  pi=24'b000000010001100100011101;
#1 $display("%b", po);
# 1  pi=24'b110011111110110001001001;
#1 $display("%b", po);
# 1  pi=24'b100010111000111001011110;
#1 $display("%b", po);
# 1  pi=24'b111011111110110000011000;
#1 $display("%b", po);
# 1  pi=24'b101001101100000010110111;
#1 $display("%b", po);
# 1  pi=24'b111100100001000001111011;
#1 $display("%b", po);
# 1  pi=24'b011111001000010011001110;
#1 $display("%b", po);
# 1  pi=24'b000001111111010011001101;
#1 $display("%b", po);
# 1  pi=24'b001010011010101010101110;
#1 $display("%b", po);
# 1  pi=24'b111001111010111001011101;
#1 $display("%b", po);
# 1  pi=24'b011011001101100001111111;
#1 $display("%b", po);
# 1  pi=24'b010001010101010011110010;
#1 $display("%b", po);
# 1  pi=24'b111110110001110110101000;
#1 $display("%b", po);
# 1  pi=24'b111010110111111010001110;
#1 $display("%b", po);
# 1  pi=24'b011110110001101000001110;
#1 $display("%b", po);
# 1  pi=24'b111010110101101000001101;
#1 $display("%b", po);
# 1  pi=24'b110111111000101111101100;
#1 $display("%b", po);
# 1  pi=24'b101010001001011011001100;
#1 $display("%b", po);
# 1  pi=24'b110010100110001101111110;
#1 $display("%b", po);
# 1  pi=24'b110011110100100110101110;
#1 $display("%b", po);
# 1  pi=24'b110011000111001100111100;
#1 $display("%b", po);
# 1  pi=24'b111110010100110111101111;
#1 $display("%b", po);
# 1  pi=24'b011000111010001000011011;
#1 $display("%b", po);
# 1  pi=24'b010001110100000111101111;
#1 $display("%b", po);
# 1  pi=24'b111001101011101001000011;
#1 $display("%b", po);
# 1  pi=24'b001011001101110101101011;
#1 $display("%b", po);
# 1  pi=24'b010010001001000111011000;
#1 $display("%b", po);
# 1  pi=24'b110001101010011100001110;
#1 $display("%b", po);
# 1  pi=24'b001110000110001111100010;
#1 $display("%b", po);
# 1  pi=24'b010000110101110001011011;
#1 $display("%b", po);
# 1  pi=24'b011011110100110000000111;
#1 $display("%b", po);
# 1  pi=24'b001100011001100101010111;
#1 $display("%b", po);
# 1  pi=24'b101100001111101011000110;
#1 $display("%b", po);
# 1  pi=24'b000011110011111110101110;
#1 $display("%b", po);
# 1  pi=24'b010011001110000100011100;
#1 $display("%b", po);
# 1  pi=24'b100110000000101000111101;
#1 $display("%b", po);
# 1  pi=24'b011111110100010101011110;
#1 $display("%b", po);
# 1  pi=24'b111111100111111111010101;
#1 $display("%b", po);
# 1  pi=24'b001101111110111110101110;
#1 $display("%b", po);
# 1  pi=24'b001110111100101101011000;
#1 $display("%b", po);
# 1  pi=24'b000011010010100101000010;
#1 $display("%b", po);
# 1  pi=24'b001010100110101010101100;
#1 $display("%b", po);
# 1  pi=24'b001101011101011100011000;
#1 $display("%b", po);
# 1  pi=24'b111010110101100001000000;
#1 $display("%b", po);
# 1  pi=24'b110011011000100110000001;
#1 $display("%b", po);
# 1  pi=24'b100001001000000101010100;
#1 $display("%b", po);
# 1  pi=24'b111000101100001110101010;
#1 $display("%b", po);
# 1  pi=24'b110110011100010101110101;
#1 $display("%b", po);
# 1  pi=24'b001001011000010000000111;
#1 $display("%b", po);
# 1  pi=24'b111111110001110000000110;
#1 $display("%b", po);
# 1  pi=24'b101100101111000010011110;
#1 $display("%b", po);
# 1  pi=24'b110100111100111111011101;
#1 $display("%b", po);
# 1  pi=24'b100101111111001101000100;
#1 $display("%b", po);
# 1  pi=24'b011000000110011001110100;
#1 $display("%b", po);
# 1  pi=24'b011001111000100110000101;
#1 $display("%b", po);
# 1  pi=24'b101110101010001100010110;
#1 $display("%b", po);
# 1  pi=24'b101110011111110000110010;
#1 $display("%b", po);
# 1  pi=24'b100000001001100000100101;
#1 $display("%b", po);
# 1  pi=24'b001011011001000000011101;
#1 $display("%b", po);
# 1  pi=24'b000111001110111100010001;
#1 $display("%b", po);
# 1  pi=24'b111010100101001101010010;
#1 $display("%b", po);
# 1  pi=24'b001100001010001000010001;
#1 $display("%b", po);
# 1  pi=24'b011011011000011011010111;
#1 $display("%b", po);
# 1  pi=24'b111110000100001001011111;
#1 $display("%b", po);
# 1  pi=24'b011100010110111001111000;
#1 $display("%b", po);
# 1  pi=24'b001100001100010001011111;
#1 $display("%b", po);
# 1  pi=24'b110010011111101111010011;
#1 $display("%b", po);
# 1  pi=24'b001110100100011111000000;
#1 $display("%b", po);
# 1  pi=24'b110001010001110001110110;
#1 $display("%b", po);
# 1  pi=24'b010011100000010101101111;
#1 $display("%b", po);
# 1  pi=24'b011000110110111000111010;
#1 $display("%b", po);
# 1  pi=24'b011010101001110100010010;
#1 $display("%b", po);
# 1  pi=24'b000101110001110101110111;
#1 $display("%b", po);
# 1  pi=24'b110000001000010001000111;
#1 $display("%b", po);
# 1  pi=24'b111100110110101110110011;
#1 $display("%b", po);
# 1  pi=24'b111001011110010101101110;
#1 $display("%b", po);
# 1  pi=24'b100101110111111011001001;
#1 $display("%b", po);
# 1  pi=24'b110010101000100101000001;
#1 $display("%b", po);
# 1  pi=24'b011011101010110010100111;
#1 $display("%b", po);
# 1  pi=24'b111111100010000011001011;
#1 $display("%b", po);
# 1  pi=24'b000110100101111101011100;
#1 $display("%b", po);
# 1  pi=24'b011100101001100100101010;
#1 $display("%b", po);
# 1  pi=24'b011100111011001110100001;
#1 $display("%b", po);
# 1  pi=24'b110110010101100111010100;
#1 $display("%b", po);
# 1  pi=24'b000001100111101110101000;
#1 $display("%b", po);
# 1  pi=24'b001011001110000111111011;
#1 $display("%b", po);
# 1  pi=24'b000010101011001111110101;
#1 $display("%b", po);
# 1  pi=24'b011111110111110010010011;
#1 $display("%b", po);
# 1  pi=24'b001001110110011010101000;
#1 $display("%b", po);
# 1  pi=24'b001010010101100011100100;
#1 $display("%b", po);
# 1  pi=24'b000001000011110111000111;
#1 $display("%b", po);
# 1  pi=24'b110010011000000110110111;
#1 $display("%b", po);
# 1  pi=24'b111001110101111111011010;
#1 $display("%b", po);
# 1  pi=24'b011000010101001110011011;
#1 $display("%b", po);
# 1  pi=24'b110111111110100010011000;
#1 $display("%b", po);
# 1  pi=24'b111110110100111110001010;
#1 $display("%b", po);
# 1  pi=24'b100011100101111111101110;
#1 $display("%b", po);
# 1  pi=24'b101111001111000010111000;
#1 $display("%b", po);
# 1  pi=24'b110111010010100100101101;
#1 $display("%b", po);
# 1  pi=24'b110110001010001011001001;
#1 $display("%b", po);
# 1  pi=24'b000110001111111101000001;
#1 $display("%b", po);
# 1  pi=24'b101101101010110110001101;
#1 $display("%b", po);
# 1  pi=24'b110011001110010000010000;
#1 $display("%b", po);
# 1  pi=24'b111111000101001001100001;
#1 $display("%b", po);
# 1  pi=24'b100101011111001110111001;
#1 $display("%b", po);
# 1  pi=24'b100001000001101010011100;
#1 $display("%b", po);
# 1  pi=24'b001110110011101010101010;
#1 $display("%b", po);
# 1  pi=24'b011110111000100111000001;
#1 $display("%b", po);
# 1  pi=24'b100101110000101001101011;
#1 $display("%b", po);
# 1  pi=24'b111011011011101110110000;
#1 $display("%b", po);
# 1  pi=24'b101011000111110001110101;
#1 $display("%b", po);
# 1  pi=24'b011000111100110010100001;
#1 $display("%b", po);
# 1  pi=24'b000111011101000111100010;
#1 $display("%b", po);
# 1  pi=24'b000100101001101000001011;
#1 $display("%b", po);
# 1  pi=24'b001110111011011100011011;
#1 $display("%b", po);
# 1  pi=24'b110110110011010000010001;
#1 $display("%b", po);
# 1  pi=24'b011011111001111100101011;
#1 $display("%b", po);
# 1  pi=24'b001110110010010000011011;
#1 $display("%b", po);
# 1  pi=24'b110011101011001110101000;
#1 $display("%b", po);
# 1  pi=24'b000110100010000110000111;
#1 $display("%b", po);
# 1  pi=24'b001110111011111011100110;
#1 $display("%b", po);
# 1  pi=24'b101110000100101000011100;
#1 $display("%b", po);
# 1  pi=24'b010101111010101011110000;
#1 $display("%b", po);
# 1  pi=24'b010100000010111010000000;
#1 $display("%b", po);
# 1  pi=24'b101001100000110100010111;
#1 $display("%b", po);
# 1  pi=24'b010000001010100011110011;
#1 $display("%b", po);
# 1  pi=24'b011011000011110111110001;
#1 $display("%b", po);
# 1  pi=24'b100111111000001010100101;
#1 $display("%b", po);
# 1  pi=24'b011111000101000111000101;
#1 $display("%b", po);
# 1  pi=24'b011100011010111000000011;
#1 $display("%b", po);
# 1  pi=24'b000110011100000100111011;
#1 $display("%b", po);
# 1  pi=24'b011110000011101010000001;
#1 $display("%b", po);
# 1  pi=24'b101000110100000010100000;
#1 $display("%b", po);
# 1  pi=24'b100011100111000100011110;
#1 $display("%b", po);
# 1  pi=24'b011011111010100001001001;
#1 $display("%b", po);
# 1  pi=24'b110010100001001011010111;
#1 $display("%b", po);
# 1  pi=24'b001011011111010010100001;
#1 $display("%b", po);
# 1  pi=24'b010101011100110111101110;
#1 $display("%b", po);
# 1  pi=24'b000101101111011110100100;
#1 $display("%b", po);
# 1  pi=24'b001111001100110001100000;
#1 $display("%b", po);
# 1  pi=24'b001011011100110011101001;
#1 $display("%b", po);
# 1  pi=24'b010101110010001000100011;
#1 $display("%b", po);
# 1  pi=24'b101001010001110010011000;
#1 $display("%b", po);
# 1  pi=24'b011111100011011010000100;
#1 $display("%b", po);
# 1  pi=24'b111110110010110100001000;
#1 $display("%b", po);
# 1  pi=24'b001001001000111000110011;
#1 $display("%b", po);
# 1  pi=24'b011110110111111000100010;
#1 $display("%b", po);
# 1  pi=24'b110001011001110110011010;
#1 $display("%b", po);
# 1  pi=24'b100011111100001100110000;
#1 $display("%b", po);
# 1  pi=24'b101010101000001000011010;
#1 $display("%b", po);
# 1  pi=24'b100110000110100111000110;
#1 $display("%b", po);
# 1  pi=24'b110001011111100110010100;
#1 $display("%b", po);
# 1  pi=24'b110010011111001110100011;
#1 $display("%b", po);
# 1  pi=24'b101011000001010100001000;
#1 $display("%b", po);
# 1  pi=24'b000000110000100001000001;
#1 $display("%b", po);
# 1  pi=24'b001000000111000011010101;
#1 $display("%b", po);
# 1  pi=24'b000110100100011010111010;
#1 $display("%b", po);
# 1  pi=24'b110100000110101010101011;
#1 $display("%b", po);
# 1  pi=24'b101101101010101110001001;
#1 $display("%b", po);
# 1  pi=24'b011100010011111111000001;
#1 $display("%b", po);
# 1  pi=24'b001100000010101100001101;
#1 $display("%b", po);
# 1  pi=24'b110111000011100001111110;
#1 $display("%b", po);
# 1  pi=24'b011110111110110000100111;
#1 $display("%b", po);
# 1  pi=24'b111101110000011100100001;
#1 $display("%b", po);
# 1  pi=24'b101111111010111011001111;
#1 $display("%b", po);
# 1  pi=24'b111100001110110111110101;
#1 $display("%b", po);
# 1  pi=24'b110110010001100000101000;
#1 $display("%b", po);
# 1  pi=24'b110001010000001011001010;
#1 $display("%b", po);
# 1  pi=24'b110001011110101111000001;
#1 $display("%b", po);
# 1  pi=24'b101100111101010101111101;
#1 $display("%b", po);
# 1  pi=24'b000000110010110100001110;
#1 $display("%b", po);
# 1  pi=24'b111010010001110101100010;
#1 $display("%b", po);
# 1  pi=24'b110110100001101000101001;
#1 $display("%b", po);
# 1  pi=24'b001100101100100101010110;
#1 $display("%b", po);
# 1  pi=24'b100110010001110110100101;
#1 $display("%b", po);
# 1  pi=24'b111100001111000101110110;
#1 $display("%b", po);
# 1  pi=24'b000100110101101001101111;
#1 $display("%b", po);
# 1  pi=24'b011000011110001111000110;
#1 $display("%b", po);
# 1  pi=24'b101101100010100110101111;
#1 $display("%b", po);
# 1  pi=24'b001110111110001110101111;
#1 $display("%b", po);
# 1  pi=24'b101010101111000110111111;
#1 $display("%b", po);
# 1  pi=24'b000101001101100111110000;
#1 $display("%b", po);
# 1  pi=24'b111011101110111000100110;
#1 $display("%b", po);
# 1  pi=24'b101011110101010010001111;
#1 $display("%b", po);
# 1  pi=24'b001000111001110001001011;
#1 $display("%b", po);
# 1  pi=24'b100111001101100010000110;
#1 $display("%b", po);
# 1  pi=24'b110111010111101001000110;
#1 $display("%b", po);
# 1  pi=24'b010110011011011011111000;
#1 $display("%b", po);
# 1  pi=24'b111000001101001010011011;
#1 $display("%b", po);
# 1  pi=24'b001101010000100000100110;
#1 $display("%b", po);
# 1  pi=24'b011010110110101100010101;
#1 $display("%b", po);
# 1  pi=24'b001101111011100100000101;
#1 $display("%b", po);
# 1  pi=24'b000111100010000000110111;
#1 $display("%b", po);
# 1  pi=24'b010000011101111100100011;
#1 $display("%b", po);
# 1  pi=24'b001101011011001101111100;
#1 $display("%b", po);
# 1  pi=24'b010010110111111101011101;
#1 $display("%b", po);
# 1  pi=24'b101000101101011000011001;
#1 $display("%b", po);
# 1  pi=24'b010001011111101111001001;
#1 $display("%b", po);
# 1  pi=24'b101110101010100101000110;
#1 $display("%b", po);
# 1  pi=24'b010101111110011100001100;
#1 $display("%b", po);
# 1  pi=24'b100111011000001001101000;
#1 $display("%b", po);
# 1  pi=24'b111110010110000100000001;
#1 $display("%b", po);
# 1  pi=24'b000100110001000110110101;
#1 $display("%b", po);
# 1  pi=24'b011011111000000110111011;
#1 $display("%b", po);
# 1  pi=24'b000001111101011110101000;
#1 $display("%b", po);
# 1  pi=24'b010111001101000000100001;
#1 $display("%b", po);
# 1  pi=24'b100110101011101000100011;
#1 $display("%b", po);
# 1  pi=24'b110101000011001100101001;
#1 $display("%b", po);
# 1  pi=24'b101010011101010100000110;
#1 $display("%b", po);
# 1  pi=24'b011110001111011011110011;
#1 $display("%b", po);
# 1  pi=24'b110011010010010001011100;
#1 $display("%b", po);
# 1  pi=24'b010101111110100001110001;
#1 $display("%b", po);
# 1  pi=24'b000110101001000001000001;
#1 $display("%b", po);
# 1  pi=24'b101011011011000100011111;
#1 $display("%b", po);
# 1  pi=24'b011101000100110001111101;
#1 $display("%b", po);
# 1  pi=24'b000111110101010011000110;
#1 $display("%b", po);
# 1  pi=24'b101110101000101101101111;
#1 $display("%b", po);
# 1  pi=24'b110101011100011011101101;
#1 $display("%b", po);
# 1  pi=24'b111011011110111001101100;
#1 $display("%b", po);
# 1  pi=24'b011111001010000010110011;
#1 $display("%b", po);
# 1  pi=24'b111110000010001100110100;
#1 $display("%b", po);
# 1  pi=24'b010000100000101110001110;
#1 $display("%b", po);
# 1  pi=24'b000110100010110110110100;
#1 $display("%b", po);
# 1  pi=24'b100000011011010000000010;
#1 $display("%b", po);
# 1  pi=24'b011001100101001100000111;
#1 $display("%b", po);
# 1  pi=24'b110101101000000001101111;
#1 $display("%b", po);
# 1  pi=24'b001101010001110001001110;
#1 $display("%b", po);
# 1  pi=24'b000000011110000110000001;
#1 $display("%b", po);
# 1  pi=24'b110110101010111111001111;
#1 $display("%b", po);
# 1  pi=24'b000100001011110001110000;
#1 $display("%b", po);
# 1  pi=24'b011110010011100110010101;
#1 $display("%b", po);
# 1  pi=24'b100111011011011000111010;
#1 $display("%b", po);
# 1  pi=24'b000110101010110110000110;
#1 $display("%b", po);
# 1  pi=24'b110101111110111010011100;
#1 $display("%b", po);
# 1  pi=24'b110011110001010101001101;
#1 $display("%b", po);
# 1  pi=24'b001111001000100111111111;
#1 $display("%b", po);
# 1  pi=24'b100011001110101110111100;
#1 $display("%b", po);
# 1  pi=24'b100011101010011011100111;
#1 $display("%b", po);
# 1  pi=24'b101010010011001011010000;
#1 $display("%b", po);
# 1  pi=24'b010011101110100010001011;
#1 $display("%b", po);
# 1  pi=24'b101100101110110101110111;
#1 $display("%b", po);
# 1  pi=24'b110001010011100010101101;
#1 $display("%b", po);
# 1  pi=24'b110100001101000010010111;
#1 $display("%b", po);
# 1  pi=24'b011010110111101111010010;
#1 $display("%b", po);
# 1  pi=24'b001111011100010000000011;
#1 $display("%b", po);
# 1  pi=24'b100101010111101011001101;
#1 $display("%b", po);
# 1  pi=24'b100110100110101001101010;
#1 $display("%b", po);
# 1  pi=24'b101100011001110011111110;
#1 $display("%b", po);
# 1  pi=24'b010100111111111000111111;
#1 $display("%b", po);
# 1  pi=24'b101111111010110110000100;
#1 $display("%b", po);
# 1  pi=24'b110010011000101001011101;
#1 $display("%b", po);
# 1  pi=24'b000011011100100001000000;
#1 $display("%b", po);
# 1  pi=24'b001001001111111011000100;
#1 $display("%b", po);
# 1  pi=24'b000111101100010100011011;
#1 $display("%b", po);
# 1  pi=24'b100011010000011111100010;
#1 $display("%b", po);
# 1  pi=24'b011111011101110110110000;
#1 $display("%b", po);
# 1  pi=24'b010001010000011100001100;
#1 $display("%b", po);
# 1  pi=24'b100110011010010001001000;
#1 $display("%b", po);
# 1  pi=24'b000100101011101100100001;
#1 $display("%b", po);
# 1  pi=24'b011001010011010111111100;
#1 $display("%b", po);
# 1  pi=24'b111011101110000101011100;
#1 $display("%b", po);
# 1  pi=24'b000000000001010011100101;
#1 $display("%b", po);
# 1  pi=24'b011000110010001110110100;
#1 $display("%b", po);
# 1  pi=24'b011000101100110111011111;
#1 $display("%b", po);
# 1  pi=24'b000001011111001101111101;
#1 $display("%b", po);
# 1  pi=24'b000010011011111110110101;
#1 $display("%b", po);
# 1  pi=24'b011110111011110000110011;
#1 $display("%b", po);
# 1  pi=24'b111111111001000011011101;
#1 $display("%b", po);
# 1  pi=24'b101000011000001100000100;
#1 $display("%b", po);
# 1  pi=24'b000110100100000000100110;
#1 $display("%b", po);
# 1  pi=24'b010000000000010101101001;
#1 $display("%b", po);
# 1  pi=24'b001010111001110101011011;
#1 $display("%b", po);
# 1  pi=24'b011010001001111000001101;
#1 $display("%b", po);
# 1  pi=24'b101100010100111100010000;
#1 $display("%b", po);
# 1  pi=24'b010010110000101001011001;
#1 $display("%b", po);
# 1  pi=24'b001110010100101100111111;
#1 $display("%b", po);
# 1  pi=24'b101100010000010001110100;
#1 $display("%b", po);
# 1  pi=24'b101110111101001100000110;
#1 $display("%b", po);
# 1  pi=24'b011110111110110110111011;
#1 $display("%b", po);
# 1  pi=24'b110111101110011000101111;
#1 $display("%b", po);
# 1  pi=24'b111011011100000101011010;
#1 $display("%b", po);
# 1  pi=24'b011000011111101001100000;
#1 $display("%b", po);
# 1  pi=24'b010101010001000010111000;
#1 $display("%b", po);
# 1  pi=24'b011100111110010001001111;
#1 $display("%b", po);
# 1  pi=24'b010001001010010110001111;
#1 $display("%b", po);
# 1  pi=24'b010000010000010111011101;
#1 $display("%b", po);
# 1  pi=24'b100100011101100110101111;
#1 $display("%b", po);
# 1  pi=24'b100000100010000101010111;
#1 $display("%b", po);
# 1  pi=24'b001110100100111010100101;
#1 $display("%b", po);
# 1  pi=24'b000100101010111100100110;
#1 $display("%b", po);
# 1  pi=24'b111100000011011010100111;
#1 $display("%b", po);
# 1  pi=24'b111001000001001110000111;
#1 $display("%b", po);
# 1  pi=24'b110011101110100010111011;
#1 $display("%b", po);
# 1  pi=24'b001010011101010111011000;
#1 $display("%b", po);
# 1  pi=24'b010010110001000001100100;
#1 $display("%b", po);
# 1  pi=24'b001010100000011111000111;
#1 $display("%b", po);
# 1  pi=24'b000110011010011010011110;
#1 $display("%b", po);
# 1  pi=24'b111100010001001011001010;
#1 $display("%b", po);
# 1  pi=24'b011101001100000100001001;
#1 $display("%b", po);
# 1  pi=24'b110101111001101110101000;
#1 $display("%b", po);
# 1  pi=24'b010000001011110011010000;
#1 $display("%b", po);
# 1  pi=24'b110110111110101101111000;
#1 $display("%b", po);
# 1  pi=24'b101001011010000101000111;
#1 $display("%b", po);
# 1  pi=24'b011000001100110000111110;
#1 $display("%b", po);
# 1  pi=24'b010100110101110100110110;
#1 $display("%b", po);
# 1  pi=24'b000101001100000001000101;
#1 $display("%b", po);
# 1  pi=24'b011111010010100101011111;
#1 $display("%b", po);
# 1  pi=24'b011110010011101111100111;
#1 $display("%b", po);
# 1  pi=24'b110010000100000100111001;
#1 $display("%b", po);
# 1  pi=24'b011110100010100011010110;
#1 $display("%b", po);
# 1  pi=24'b011101101111011011010100;
#1 $display("%b", po);
# 1  pi=24'b101110000110000011000000;
#1 $display("%b", po);
# 1  pi=24'b111101010011000101010001;
#1 $display("%b", po);
# 1  pi=24'b011010000111001011111101;
#1 $display("%b", po);
# 1  pi=24'b101101011100101000100000;
#1 $display("%b", po);
# 1  pi=24'b001101101100111100100100;
#1 $display("%b", po);
# 1  pi=24'b111010110011101101010110;
#1 $display("%b", po);
# 1  pi=24'b001100100010100100010111;
#1 $display("%b", po);
# 1  pi=24'b011100111010100010010011;
#1 $display("%b", po);
# 1  pi=24'b100001111101101000000110;
#1 $display("%b", po);
# 1  pi=24'b011101100101001101010010;
#1 $display("%b", po);
# 1  pi=24'b100101010100101111001000;
#1 $display("%b", po);
# 1  pi=24'b101100111011110110110010;
#1 $display("%b", po);
# 1  pi=24'b100111011111000011011110;
#1 $display("%b", po);
# 1  pi=24'b010110110001101011111000;
#1 $display("%b", po);
# 1  pi=24'b001111001001001011111100;
#1 $display("%b", po);
# 1  pi=24'b101011101000010001000101;
#1 $display("%b", po);
# 1  pi=24'b101010111100010000010001;
#1 $display("%b", po);
# 1  pi=24'b110111110010000111110111;
#1 $display("%b", po);
# 1  pi=24'b000010110010111111010011;
#1 $display("%b", po);
# 1  pi=24'b010101111001000101001110;
#1 $display("%b", po);
# 1  pi=24'b101101110111100000111011;
#1 $display("%b", po);
# 1  pi=24'b100111010010110100000110;
#1 $display("%b", po);
# 1  pi=24'b011100110000111101101100;
#1 $display("%b", po);
# 1  pi=24'b001100001011011011111010;
#1 $display("%b", po);
# 1  pi=24'b110110011000000110100111;
#1 $display("%b", po);
# 1  pi=24'b111001100111100010100111;
#1 $display("%b", po);
# 1  pi=24'b000011001111010011100010;
#1 $display("%b", po);
# 1  pi=24'b110010010001011111110111;
#1 $display("%b", po);
# 1  pi=24'b111010110011011000110001;
#1 $display("%b", po);
# 1  pi=24'b111100111111001011110000;
#1 $display("%b", po);
# 1  pi=24'b110111110101111100110111;
#1 $display("%b", po);
# 1  pi=24'b001011101100011101110000;
#1 $display("%b", po);
# 1  pi=24'b011111010110010110011000;
#1 $display("%b", po);
# 1  pi=24'b110011110000100011110010;
#1 $display("%b", po);
# 1  pi=24'b010101110100001110110011;
#1 $display("%b", po);
# 1  pi=24'b011000111101001110101101;
#1 $display("%b", po);
# 1  pi=24'b111111000111011111000110;
#1 $display("%b", po);
# 1  pi=24'b011110011101010101101101;
#1 $display("%b", po);
# 1  pi=24'b010001000000000111000101;
#1 $display("%b", po);
# 1  pi=24'b111111110111010001111011;
#1 $display("%b", po);
# 1  pi=24'b101110011011110110111000;
#1 $display("%b", po);
# 1  pi=24'b011100010011101000001111;
#1 $display("%b", po);
# 1  pi=24'b001010000111010001101011;
#1 $display("%b", po);
# 1  pi=24'b010101000011101100010010;
#1 $display("%b", po);
# 1  pi=24'b011101101001100000011101;
#1 $display("%b", po);
# 1  pi=24'b011111101011011001000001;
#1 $display("%b", po);
# 1  pi=24'b001101100110010110011101;
#1 $display("%b", po);
# 1  pi=24'b111101000110100001011011;
#1 $display("%b", po);
# 1  pi=24'b011011001001010101010000;
#1 $display("%b", po);
# 1  pi=24'b000001001011110001100111;
#1 $display("%b", po);
# 1  pi=24'b101111110101101000111001;
#1 $display("%b", po);
# 1  pi=24'b011110100000110111100101;
#1 $display("%b", po);
# 1  pi=24'b100001110110100101100000;
#1 $display("%b", po);
# 1  pi=24'b010101111000011100100010;
#1 $display("%b", po);
# 1  pi=24'b100010001110110111011111;
#1 $display("%b", po);
# 1  pi=24'b001000011111100110101101;
#1 $display("%b", po);
# 1  pi=24'b000111000111001011011101;
#1 $display("%b", po);
# 1  pi=24'b111000101100011110011111;
#1 $display("%b", po);
# 1  pi=24'b001100100110001011000100;
#1 $display("%b", po);
# 1  pi=24'b111101011001001110010111;
#1 $display("%b", po);
# 1  pi=24'b000110110001100000010011;
#1 $display("%b", po);
# 1  pi=24'b001010110110011110111000;
#1 $display("%b", po);
# 1  pi=24'b110001011001010110110110;
#1 $display("%b", po);
# 1  pi=24'b101001010101100010110100;
#1 $display("%b", po);
# 1  pi=24'b100010110100111101111000;
#1 $display("%b", po);
# 1  pi=24'b011000000100111000001101;
#1 $display("%b", po);
# 1  pi=24'b110101111010110101110000;
#1 $display("%b", po);
# 1  pi=24'b010101000001100010011000;
#1 $display("%b", po);
# 1  pi=24'b000001011111110100111100;
#1 $display("%b", po);
# 1  pi=24'b100010000010100011111010;
#1 $display("%b", po);
# 1  pi=24'b111100100111011111000100;
#1 $display("%b", po);
# 1  pi=24'b001100000110100111100100;
#1 $display("%b", po);
# 1  pi=24'b101110100100010000110011;
#1 $display("%b", po);
# 1  pi=24'b010000111111101010011111;
#1 $display("%b", po);
# 1  pi=24'b100001011011101100101000;
#1 $display("%b", po);
# 1  pi=24'b101101010010001010011100;
#1 $display("%b", po);
# 1  pi=24'b000001000111011110100101;
#1 $display("%b", po);
# 1  pi=24'b111100010100001010100010;
#1 $display("%b", po);
# 1  pi=24'b110000100101101000011111;
#1 $display("%b", po);
# 1  pi=24'b111001010110001110100100;
#1 $display("%b", po);
# 1  pi=24'b110010011011100100010101;
#1 $display("%b", po);
# 1  pi=24'b100101011110001000100100;
#1 $display("%b", po);
# 1  pi=24'b001010101001001100001100;
#1 $display("%b", po);
# 1  pi=24'b110000101100000010010111;
#1 $display("%b", po);
# 1  pi=24'b110001001010100101100001;
#1 $display("%b", po);
# 1  pi=24'b010111101011011011001110;
#1 $display("%b", po);
# 1  pi=24'b010100000010001010101110;
#1 $display("%b", po);
# 1  pi=24'b001100000100101110111011;
#1 $display("%b", po);
# 1  pi=24'b111100001110100011010011;
#1 $display("%b", po);
# 1  pi=24'b000011000100001101011011;
#1 $display("%b", po);
# 1  pi=24'b110000000011010010111000;
#1 $display("%b", po);
# 1  pi=24'b001001000111011100011010;
#1 $display("%b", po);
# 1  pi=24'b010001011010110100111011;
#1 $display("%b", po);
# 1  pi=24'b101010001011111100001011;
#1 $display("%b", po);
# 1  pi=24'b101011011100000010110001;
#1 $display("%b", po);
# 1  pi=24'b101101100101101011010101;
#1 $display("%b", po);
# 1  pi=24'b100100110001101011011011;
#1 $display("%b", po);
# 1  pi=24'b010111011101000100011001;
#1 $display("%b", po);
# 1  pi=24'b001000110001101010010101;
#1 $display("%b", po);
# 1  pi=24'b100011001010010110101011;
#1 $display("%b", po);
# 1  pi=24'b111010000100100000110100;
#1 $display("%b", po);
# 1  pi=24'b101000010100101111000011;
#1 $display("%b", po);
# 1  pi=24'b101111011010110110111111;
#1 $display("%b", po);
# 1  pi=24'b101100100000110011011110;
#1 $display("%b", po);
# 1  pi=24'b000101111000001101101011;
#1 $display("%b", po);
# 1  pi=24'b110110101001001111011101;
#1 $display("%b", po);
# 1  pi=24'b011011111010101010111001;
#1 $display("%b", po);
# 1  pi=24'b100110100000100001110001;
#1 $display("%b", po);
# 1  pi=24'b100010000010110011011001;
#1 $display("%b", po);
# 1  pi=24'b000011011111101100100111;
#1 $display("%b", po);
# 1  pi=24'b001110111101101010110101;
#1 $display("%b", po);
# 1  pi=24'b000010110001011011100010;
#1 $display("%b", po);
# 1  pi=24'b010010101111111110001110;
#1 $display("%b", po);
# 1  pi=24'b110011100001100100010101;
#1 $display("%b", po);
# 1  pi=24'b011100110000111011010000;
#1 $display("%b", po);
# 1  pi=24'b011101000011111110100100;
#1 $display("%b", po);
# 1  pi=24'b110001100111011011101100;
#1 $display("%b", po);
# 1  pi=24'b100011110101110001010000;
#1 $display("%b", po);
# 1  pi=24'b011001011001111111111000;
#1 $display("%b", po);
# 1  pi=24'b001110100011110100000101;
#1 $display("%b", po);
# 1  pi=24'b011010000111010110000000;
#1 $display("%b", po);
# 1  pi=24'b101010000110001011010100;
#1 $display("%b", po);
# 1  pi=24'b101011110100101111000111;
#1 $display("%b", po);
# 1  pi=24'b110100100000001111100100;
#1 $display("%b", po);
# 1  pi=24'b111010100011111101110010;
#1 $display("%b", po);
# 1  pi=24'b111001100110100000111010;
#1 $display("%b", po);
# 1  pi=24'b110001010111001100000111;
#1 $display("%b", po);
# 1  pi=24'b011101001101010001010001;
#1 $display("%b", po);
# 1  pi=24'b111010010011110011010100;
#1 $display("%b", po);
# 1  pi=24'b001100111000111111001001;
#1 $display("%b", po);
# 1  pi=24'b011000110000010100111111;
#1 $display("%b", po);
# 1  pi=24'b001100110000100000010010;
#1 $display("%b", po);
# 1  pi=24'b101111001001111100001000;
#1 $display("%b", po);
# 1  pi=24'b101011111101111000010011;
#1 $display("%b", po);
# 1  pi=24'b111010010111110010100101;
#1 $display("%b", po);
# 1  pi=24'b001000010101100000011101;
#1 $display("%b", po);
# 1  pi=24'b011010010011110110001010;
#1 $display("%b", po);
# 1  pi=24'b111100110111001000010010;
#1 $display("%b", po);
# 1  pi=24'b101100100001001111101101;
#1 $display("%b", po);
# 1  pi=24'b010100101101001000111011;
#1 $display("%b", po);
# 1  pi=24'b011110000011100000110100;
#1 $display("%b", po);
# 1  pi=24'b011000101101100100101110;
#1 $display("%b", po);
# 1  pi=24'b100100100100000011101011;
#1 $display("%b", po);
# 1  pi=24'b001110010001001101111111;
#1 $display("%b", po);
# 1  pi=24'b001100111010001011101110;
#1 $display("%b", po);
# 1  pi=24'b101111101100011110100101;
#1 $display("%b", po);
# 1  pi=24'b111001101111010001011011;
#1 $display("%b", po);
# 1  pi=24'b001001110100011110101111;
#1 $display("%b", po);
# 1  pi=24'b110100010110110010100110;
#1 $display("%b", po);
# 1  pi=24'b010101011101000100100000;
#1 $display("%b", po);
# 1  pi=24'b011110011001011011001111;
#1 $display("%b", po);
# 1  pi=24'b000101010010000000111001;
#1 $display("%b", po);
# 1  pi=24'b111011010110010000001011;
#1 $display("%b", po);
# 1  pi=24'b110100001101101100010111;
#1 $display("%b", po);
# 1  pi=24'b110110010010011111010000;
#1 $display("%b", po);
# 1  pi=24'b111111001001100111110111;
#1 $display("%b", po);
# 1  pi=24'b110101110010111100011010;
#1 $display("%b", po);
# 1  pi=24'b001101111110100100011001;
#1 $display("%b", po);
# 1  pi=24'b100011101001110011110010;
#1 $display("%b", po);
# 1  pi=24'b000000101011111110001001;
#1 $display("%b", po);
# 1  pi=24'b100011111000110101100010;
#1 $display("%b", po);
# 1  pi=24'b000011000111001010110001;
#1 $display("%b", po);
# 1  pi=24'b010111001011100010110110;
#1 $display("%b", po);
# 1  pi=24'b101001101000100011111010;
#1 $display("%b", po);
# 1  pi=24'b010100100111010110101101;
#1 $display("%b", po);
# 1  pi=24'b100110000010001000100101;
#1 $display("%b", po);
# 1  pi=24'b101110111001001110000100;
#1 $display("%b", po);
# 1  pi=24'b001110111101100111011100;
#1 $display("%b", po);
# 1  pi=24'b111110100001110111010000;
#1 $display("%b", po);
# 1  pi=24'b010011100101110101110110;
#1 $display("%b", po);
# 1  pi=24'b011001010010011111101100;
#1 $display("%b", po);
# 1  pi=24'b011110001001000111001011;
#1 $display("%b", po);
# 1  pi=24'b111100001001000001001100;
#1 $display("%b", po);
# 1  pi=24'b101100110011000100111001;
#1 $display("%b", po);
# 1  pi=24'b111000000001101100001010;
#1 $display("%b", po);
# 1  pi=24'b011111100010011011111110;
#1 $display("%b", po);
# 1  pi=24'b000100110110011001000010;
#1 $display("%b", po);
# 1  pi=24'b110110101000101010110110;
#1 $display("%b", po);
# 1  pi=24'b001110110010011000110111;
#1 $display("%b", po);
# 1  pi=24'b000011110001011110101111;
#1 $display("%b", po);
# 1  pi=24'b000110110010010110011000;
#1 $display("%b", po);
# 1  pi=24'b000111101101001101110010;
#1 $display("%b", po);
# 1  pi=24'b101110011001110101010101;
#1 $display("%b", po);
# 1  pi=24'b000111001010001110011110;
#1 $display("%b", po);
# 1  pi=24'b110001110000101100001110;
#1 $display("%b", po);
# 1  pi=24'b010110011110101000111100;
#1 $display("%b", po);
# 1  pi=24'b010111001000111111110010;
#1 $display("%b", po);
# 1  pi=24'b101100000111100001000000;
#1 $display("%b", po);
# 1  pi=24'b011011000101000010001111;
#1 $display("%b", po);
# 1  pi=24'b000000010101101100000110;
#1 $display("%b", po);
# 1  pi=24'b001010001011101100001001;
#1 $display("%b", po);
# 1  pi=24'b000110000111110111110001;
#1 $display("%b", po);
# 1  pi=24'b111100100101101001110000;
#1 $display("%b", po);
# 1  pi=24'b100101111110000001001010;
#1 $display("%b", po);
# 1  pi=24'b100000110010101001001001;
#1 $display("%b", po);
# 1  pi=24'b010100010000000001001011;
#1 $display("%b", po);
# 1  pi=24'b001100011001000100111011;
#1 $display("%b", po);
# 1  pi=24'b111111101001001111110000;
#1 $display("%b", po);
# 1  pi=24'b100110100000100010110100;
#1 $display("%b", po);
# 1  pi=24'b001101000001011010101010;
#1 $display("%b", po);
# 1  pi=24'b001111111000110001100111;
#1 $display("%b", po);
# 1  pi=24'b000011011000000111101010;
#1 $display("%b", po);
# 1  pi=24'b101000000011010001101001;
#1 $display("%b", po);
# 1  pi=24'b110011100110011001100001;
#1 $display("%b", po);
# 1  pi=24'b010100100010000100011011;
#1 $display("%b", po);
# 1  pi=24'b000011001001100011011110;
#1 $display("%b", po);
# 1  pi=24'b101010100101000000000000;
#1 $display("%b", po);
# 1  pi=24'b101111010000010100010001;
#1 $display("%b", po);
# 1  pi=24'b100110000000101100110001;
#1 $display("%b", po);
# 1  pi=24'b011111010100100000010001;
#1 $display("%b", po);
# 1  pi=24'b111101011101111100111101;
#1 $display("%b", po);
# 1  pi=24'b010000110011100101101100;
#1 $display("%b", po);
# 1  pi=24'b000011010000001100011101;
#1 $display("%b", po);
# 1  pi=24'b111110011000011010000001;
#1 $display("%b", po);
# 1  pi=24'b000110111110010111001101;
#1 $display("%b", po);
# 1  pi=24'b010100001011011110110011;
#1 $display("%b", po);
# 1  pi=24'b001010100101010000001010;
#1 $display("%b", po);
# 1  pi=24'b110100011001101101101101;
#1 $display("%b", po);
# 1  pi=24'b110011001100000010000101;
#1 $display("%b", po);
# 1  pi=24'b110001111001010010011110;
#1 $display("%b", po);
# 1  pi=24'b000101111011110000011010;
#1 $display("%b", po);
# 1  pi=24'b010001011111001110001000;
#1 $display("%b", po);
# 1  pi=24'b001111101101000111100100;
#1 $display("%b", po);
# 1  pi=24'b100101101001110110100000;
#1 $display("%b", po);
# 1  pi=24'b010111110100111011000111;
#1 $display("%b", po);
# 1  pi=24'b100000110011011100000010;
#1 $display("%b", po);
# 1  pi=24'b100001001100111010010100;
#1 $display("%b", po);
# 1  pi=24'b011010100101110111010110;
#1 $display("%b", po);
# 1  pi=24'b111010010111100100000001;
#1 $display("%b", po);
# 1  pi=24'b001001100011010110011011;
#1 $display("%b", po);
# 1  pi=24'b101010100010000010001011;
#1 $display("%b", po);
# 1  pi=24'b111110011001101100111001;
#1 $display("%b", po);
# 1  pi=24'b101100000000111111000110;
#1 $display("%b", po);
# 1  pi=24'b000001101001011101110110;
#1 $display("%b", po);
# 1  pi=24'b111010101100101111101100;
#1 $display("%b", po);
# 1  pi=24'b110000000111111100111000;
#1 $display("%b", po);
# 1  pi=24'b010111011111001111110001;
#1 $display("%b", po);
# 1  pi=24'b001110011010111111010111;
#1 $display("%b", po);
# 1  pi=24'b110011001010000001000011;
#1 $display("%b", po);
# 1  pi=24'b000000010010011010110101;
#1 $display("%b", po);
# 1  pi=24'b100011010000100100011011;
#1 $display("%b", po);
# 1  pi=24'b011100111010000101101100;
#1 $display("%b", po);
# 1  pi=24'b000001100011100011101001;
#1 $display("%b", po);
# 1  pi=24'b111110000010010011011111;
#1 $display("%b", po);
# 1  pi=24'b011000000010101011101010;
#1 $display("%b", po);
# 1  pi=24'b001101100111100000000100;
#1 $display("%b", po);
# 1  pi=24'b111111111000110010011111;
#1 $display("%b", po);
# 1  pi=24'b101010001000010110010000;
#1 $display("%b", po);
# 1  pi=24'b001010001101110001101101;
#1 $display("%b", po);
# 1  pi=24'b100011000110010011100001;
#1 $display("%b", po);
# 1  pi=24'b000011111001111001011110;
#1 $display("%b", po);
# 1  pi=24'b010001011001010101011011;
#1 $display("%b", po);
# 1  pi=24'b011011011111001100100000;
#1 $display("%b", po);
# 1  pi=24'b101000100111110010001001;
#1 $display("%b", po);
# 1  pi=24'b000100011111010110100000;
#1 $display("%b", po);
# 1  pi=24'b110011001110100101000111;
#1 $display("%b", po);
# 1  pi=24'b101011010011000100101011;
#1 $display("%b", po);
# 1  pi=24'b001010100000010101011111;
#1 $display("%b", po);
# 1  pi=24'b001101101101111101101100;
#1 $display("%b", po);
# 1  pi=24'b100111001111011001000101;
#1 $display("%b", po);
# 1  pi=24'b001110011110111100011010;
#1 $display("%b", po);
# 1  pi=24'b100101000010101100001110;
#1 $display("%b", po);
# 1  pi=24'b110010011001011000001111;
#1 $display("%b", po);
# 1  pi=24'b101111111000000000001000;
#1 $display("%b", po);
# 1  pi=24'b110011101101001100010100;
#1 $display("%b", po);
# 1  pi=24'b101010011100011001011000;
#1 $display("%b", po);
# 1  pi=24'b000100001111001111101100;
#1 $display("%b", po);
# 1  pi=24'b101100101000111000000111;
#1 $display("%b", po);
# 1  pi=24'b111000101111001110101100;
#1 $display("%b", po);
# 1  pi=24'b000011000111011101000110;
#1 $display("%b", po);
# 1  pi=24'b100011010110001010110011;
#1 $display("%b", po);
# 1  pi=24'b001110001010000001110110;
#1 $display("%b", po);
# 1  pi=24'b111000111111000101100101;
#1 $display("%b", po);
# 1  pi=24'b001100111110111001110010;
#1 $display("%b", po);
# 1  pi=24'b011001110011000110010110;
#1 $display("%b", po);
# 1  pi=24'b001100011010100100011000;
#1 $display("%b", po);
# 1  pi=24'b100101101101010110100100;
#1 $display("%b", po);
# 1  pi=24'b000011100000111111010001;
#1 $display("%b", po);
# 1  pi=24'b110101100101001110000111;
#1 $display("%b", po);
# 1  pi=24'b111111000010001100011011;
#1 $display("%b", po);
# 1  pi=24'b000001110111100111011011;
#1 $display("%b", po);
# 1  pi=24'b001110101100111111101001;
#1 $display("%b", po);
# 1  pi=24'b111101010100011000100011;
#1 $display("%b", po);
# 1  pi=24'b010111100110101000101011;
#1 $display("%b", po);
# 1  pi=24'b010010000101100111000001;
#1 $display("%b", po);
# 1  pi=24'b001001111000111110001111;
#1 $display("%b", po);
# 1  pi=24'b101011001100000011110010;
#1 $display("%b", po);
# 1  pi=24'b000100110011000011110000;
#1 $display("%b", po);
# 1  pi=24'b010010001100010110011011;
#1 $display("%b", po);
# 1  pi=24'b110000100100100001001000;
#1 $display("%b", po);
# 1  pi=24'b101100000001010111110010;
#1 $display("%b", po);
# 1  pi=24'b011001111101011100001110;
#1 $display("%b", po);
# 1  pi=24'b001110100111100011010110;
#1 $display("%b", po);
# 1  pi=24'b100001001011001110111010;
#1 $display("%b", po);
# 1  pi=24'b001110000001100101100110;
#1 $display("%b", po);
# 1  pi=24'b111001101101110010100100;
#1 $display("%b", po);
# 1  pi=24'b000100001001100010100000;
#1 $display("%b", po);
# 1  pi=24'b110011000001001000111011;
#1 $display("%b", po);
# 1  pi=24'b011011001010000000101101;
#1 $display("%b", po);
# 1  pi=24'b101001110111011101000000;
#1 $display("%b", po);
# 1  pi=24'b010100111101001110010110;
#1 $display("%b", po);
# 1  pi=24'b010000011001011001101111;
#1 $display("%b", po);
# 1  pi=24'b101100011010001001010110;
#1 $display("%b", po);
# 1  pi=24'b010000100100000010011000;
#1 $display("%b", po);
# 1  pi=24'b000000110001011101001011;
#1 $display("%b", po);
# 1  pi=24'b110110010001110001001000;
#1 $display("%b", po);
# 1  pi=24'b011010011110010111000001;
#1 $display("%b", po);
# 1  pi=24'b100010001010000000010101;
#1 $display("%b", po);
# 1  pi=24'b100011101011100000001111;
#1 $display("%b", po);
# 1  pi=24'b100011001011101100001110;
#1 $display("%b", po);
# 1  pi=24'b000101101010010111000011;
#1 $display("%b", po);
# 1  pi=24'b111101011100101000000010;
#1 $display("%b", po);
# 1  pi=24'b100110101111011001010011;
#1 $display("%b", po);
# 1  pi=24'b101111111111110010100111;
#1 $display("%b", po);
# 1  pi=24'b010010101010000101000110;
#1 $display("%b", po);
# 1  pi=24'b010011010011000011011001;
#1 $display("%b", po);
# 1  pi=24'b111001010010100101111011;
#1 $display("%b", po);
# 1  pi=24'b001001010000101101010000;
#1 $display("%b", po);
# 1  pi=24'b010110111110000000000011;
#1 $display("%b", po);
# 1  pi=24'b101101111101001011101100;
#1 $display("%b", po);
# 1  pi=24'b100001010100110011100100;
#1 $display("%b", po);
# 1  pi=24'b100110001001001110110001;
#1 $display("%b", po);
# 1  pi=24'b110001000100001010001110;
#1 $display("%b", po);
# 1  pi=24'b101001011111000100010101;
#1 $display("%b", po);
# 1  pi=24'b011011100001011101010111;
#1 $display("%b", po);
# 1  pi=24'b011101110010001111000011;
#1 $display("%b", po);
# 1  pi=24'b110101011100100101111101;
#1 $display("%b", po);
# 1  pi=24'b001011001110110111011001;
#1 $display("%b", po);
# 1  pi=24'b100000111100100011111001;
#1 $display("%b", po);
# 1  pi=24'b010100101011110011011100;
#1 $display("%b", po);
# 1  pi=24'b011101011011000010110001;
#1 $display("%b", po);
# 1  pi=24'b000000100011010100011000;
#1 $display("%b", po);
# 1  pi=24'b111110100010011111110000;
#1 $display("%b", po);
# 1  pi=24'b000101100001110001100100;
#1 $display("%b", po);
# 1  pi=24'b111000000101100111000101;
#1 $display("%b", po);
# 1  pi=24'b001100110011101100110110;
#1 $display("%b", po);
# 1  pi=24'b011111011100111101100010;
#1 $display("%b", po);
# 1  pi=24'b011000000000110010001111;
#1 $display("%b", po);
# 1  pi=24'b110011111110111111101010;
#1 $display("%b", po);
# 1  pi=24'b010101011010100100111000;
#1 $display("%b", po);
# 1  pi=24'b010010001000111110011011;
#1 $display("%b", po);
# 1  pi=24'b001110101101010110011111;
#1 $display("%b", po);
# 1  pi=24'b110010010111101100110011;
#1 $display("%b", po);
# 1  pi=24'b000101000000101110001001;
#1 $display("%b", po);
# 1  pi=24'b111101101100111011001100;
#1 $display("%b", po);
# 1  pi=24'b101100110111100000100000;
#1 $display("%b", po);
# 1  pi=24'b000110010001101011101110;
#1 $display("%b", po);
# 1  pi=24'b000110100010110101110000;
#1 $display("%b", po);
# 1  pi=24'b110101011111111010010111;
#1 $display("%b", po);
# 1  pi=24'b010000110001001010101001;
#1 $display("%b", po);
# 1  pi=24'b101110001011000111011110;
#1 $display("%b", po);
# 1  pi=24'b000111110001001110100110;
#1 $display("%b", po);
# 1  pi=24'b010000000101101010001111;
#1 $display("%b", po);
# 1  pi=24'b011011011101010000101010;
#1 $display("%b", po);
# 1  pi=24'b010011111110000000001011;
#1 $display("%b", po);
# 1  pi=24'b001110110110101011001011;
#1 $display("%b", po);
# 1  pi=24'b101110100100100101001010;
#1 $display("%b", po);
# 1  pi=24'b011111111101100001010000;
#1 $display("%b", po);
# 1  pi=24'b101111001011100110010110;
#1 $display("%b", po);
# 1  pi=24'b011010110111111001000111;
#1 $display("%b", po);
# 1  pi=24'b110110000011111101111111;
#1 $display("%b", po);
# 1  pi=24'b010010101100111110111100;
#1 $display("%b", po);
# 1  pi=24'b011101110101011100101111;
#1 $display("%b", po);
# 1  pi=24'b010111010111100100101110;
#1 $display("%b", po);
# 1  pi=24'b011001000111110001011111;
#1 $display("%b", po);
# 1  pi=24'b101010100011111010011001;
#1 $display("%b", po);
# 1  pi=24'b000001111100101110111100;
#1 $display("%b", po);
# 1  pi=24'b111011011111001111111101;
#1 $display("%b", po);
# 1  pi=24'b110001010001001001011011;
#1 $display("%b", po);
# 1  pi=24'b010100010111011111100100;
#1 $display("%b", po);
# 1  pi=24'b101101000011111011100010;
#1 $display("%b", po);
# 1  pi=24'b110111110010100101111110;
#1 $display("%b", po);
# 1  pi=24'b101001001000010110111011;
#1 $display("%b", po);
# 1  pi=24'b100110100000010010001011;
#1 $display("%b", po);
# 1  pi=24'b011110111011101011100011;
#1 $display("%b", po);
# 1  pi=24'b000011010011101010101111;
#1 $display("%b", po);
# 1  pi=24'b011001000000111111100110;
#1 $display("%b", po);
# 1  pi=24'b010111000111010001001100;
#1 $display("%b", po);
# 1  pi=24'b011000110000101010000101;
#1 $display("%b", po);
# 1  pi=24'b111101001111000010000100;
#1 $display("%b", po);
# 1  pi=24'b001100101001001101010101;
#1 $display("%b", po);
# 1  pi=24'b011101001100001011110101;
#1 $display("%b", po);
# 1  pi=24'b100110110110010000011001;
#1 $display("%b", po);
# 1  pi=24'b111100110000110111110111;
#1 $display("%b", po);
# 1  pi=24'b111100110000011010011101;
#1 $display("%b", po);
# 1  pi=24'b100010011111000110011010;
#1 $display("%b", po);
# 1  pi=24'b000011110100100100001011;
#1 $display("%b", po);
# 1  pi=24'b011110100010111010110000;
#1 $display("%b", po);
# 1  pi=24'b011111001011101100010000;
#1 $display("%b", po);
# 1  pi=24'b100011001001000101010101;
#1 $display("%b", po);
# 1  pi=24'b001101111101110010000111;
#1 $display("%b", po);
# 1  pi=24'b001100110000100101110010;
#1 $display("%b", po);
# 1  pi=24'b110110000001010010110000;
#1 $display("%b", po);
# 1  pi=24'b011011010111100110111101;
#1 $display("%b", po);
# 1  pi=24'b011011110000100010011110;
#1 $display("%b", po);
# 1  pi=24'b100000000001100110111101;
#1 $display("%b", po);
# 1  pi=24'b100000111110010000111100;
#1 $display("%b", po);
# 1  pi=24'b011111010110011011001000;
#1 $display("%b", po);
# 1  pi=24'b101011100001001010110000;
#1 $display("%b", po);
# 1  pi=24'b101011011110001100101010;
#1 $display("%b", po);
# 1  pi=24'b100100011101100011011011;
#1 $display("%b", po);
# 1  pi=24'b010111100100111010010010;
#1 $display("%b", po);
# 1  pi=24'b110111011001110000101100;
#1 $display("%b", po);
# 1  pi=24'b110100010000001110110010;
#1 $display("%b", po);
# 1  pi=24'b100110001101101001100000;
#1 $display("%b", po);
# 1  pi=24'b000011000101000011000110;
#1 $display("%b", po);
# 1  pi=24'b000100111011110001011101;
#1 $display("%b", po);
# 1  pi=24'b000000011001000010010111;
#1 $display("%b", po);
# 1  pi=24'b010000000100011100111001;
#1 $display("%b", po);
# 1  pi=24'b010101001110101100110111;
#1 $display("%b", po);
# 1  pi=24'b010000001000110011110100;
#1 $display("%b", po);
# 1  pi=24'b011101000100111111000011;
#1 $display("%b", po);
# 1  pi=24'b111010101001110101011010;
#1 $display("%b", po);
# 1  pi=24'b001110110001001100100001;
#1 $display("%b", po);
# 1  pi=24'b101111111001010011000000;
#1 $display("%b", po);
# 1  pi=24'b010000000001111100000000;
#1 $display("%b", po);
# 1  pi=24'b110000110011010000010111;
#1 $display("%b", po);
# 1  pi=24'b010000011001010111110000;
#1 $display("%b", po);
# 1  pi=24'b011001001001010100111011;
#1 $display("%b", po);
# 1  pi=24'b001010011000001001010100;
#1 $display("%b", po);
# 1  pi=24'b010000111111010101111010;
#1 $display("%b", po);
# 1  pi=24'b010100111011000001101101;
#1 $display("%b", po);
# 1  pi=24'b101011110010011001100101;
#1 $display("%b", po);
# 1  pi=24'b010101001000000110010010;
#1 $display("%b", po);
# 1  pi=24'b110101101010111000100010;
#1 $display("%b", po);
# 1  pi=24'b010100111110100111101011;
#1 $display("%b", po);
# 1  pi=24'b111111111010001100100010;
#1 $display("%b", po);
# 1  pi=24'b011010010111000110111011;
#1 $display("%b", po);
# 1  pi=24'b001000010001110000000010;
#1 $display("%b", po);
# 1  pi=24'b111101001110011100101011;
#1 $display("%b", po);
# 1  pi=24'b010010100101001001000100;
#1 $display("%b", po);
# 1  pi=24'b000111010001000111010001;
#1 $display("%b", po);
# 1  pi=24'b100001011000011010101001;
#1 $display("%b", po);
# 1  pi=24'b100101101010010100111111;
#1 $display("%b", po);
# 1  pi=24'b101000000001010000000000;
#1 $display("%b", po);
# 1  pi=24'b001010111010010000100111;
#1 $display("%b", po);
# 1  pi=24'b111010011010101110001011;
#1 $display("%b", po);
# 1  pi=24'b111010111101110111011111;
#1 $display("%b", po);
# 1  pi=24'b000010011000111110100010;
#1 $display("%b", po);
# 1  pi=24'b010110100100110010011011;
#1 $display("%b", po);
# 1  pi=24'b111110010111111010111111;
#1 $display("%b", po);
# 1  pi=24'b100000000010001100010000;
#1 $display("%b", po);
# 1  pi=24'b100001111111000110001010;
#1 $display("%b", po);
# 1  pi=24'b111010101111001100101010;
#1 $display("%b", po);
# 1  pi=24'b101111010011100110101010;
#1 $display("%b", po);
# 1  pi=24'b110001011101011001011101;
#1 $display("%b", po);
# 1  pi=24'b001101100001010011101011;
#1 $display("%b", po);
# 1  pi=24'b010001011001110011001110;
#1 $display("%b", po);
# 1  pi=24'b100110011100110011011010;
#1 $display("%b", po);
# 1  pi=24'b111001100110110010111011;
#1 $display("%b", po);
# 1  pi=24'b111000101111000101111001;
#1 $display("%b", po);
# 1  pi=24'b011100100011100001101001;
#1 $display("%b", po);
# 1  pi=24'b001101111000000010111011;
#1 $display("%b", po);
# 1  pi=24'b011001011110111001111001;
#1 $display("%b", po);
# 1  pi=24'b110111100110010100010011;
#1 $display("%b", po);
# 1  pi=24'b001111101011000001111011;
#1 $display("%b", po);
# 1  pi=24'b111100001110010010101101;
#1 $display("%b", po);
# 1  pi=24'b101111000111101100000001;
#1 $display("%b", po);
# 1  pi=24'b111110100011011001010011;
#1 $display("%b", po);
# 1  pi=24'b000100101001110001010100;
#1 $display("%b", po);
# 1  pi=24'b010110111010010010110111;
#1 $display("%b", po);
# 1  pi=24'b111110001111000010100010;
#1 $display("%b", po);
# 1  pi=24'b110101100110010001011100;
#1 $display("%b", po);
# 1  pi=24'b100010011001010010001011;
#1 $display("%b", po);
# 1  pi=24'b101100100011111010111001;
#1 $display("%b", po);
# 1  pi=24'b101000100001101100101100;
#1 $display("%b", po);
# 1  pi=24'b110110010001110101010101;
#1 $display("%b", po);
# 1  pi=24'b111110110100110000011101;
#1 $display("%b", po);
# 1  pi=24'b010001000000111010111000;
#1 $display("%b", po);
# 1  pi=24'b001010111101010001110001;
#1 $display("%b", po);
# 1  pi=24'b001101111000101011000000;
#1 $display("%b", po);
# 1  pi=24'b111001101010111000111101;
#1 $display("%b", po);
# 1  pi=24'b110101111011101011100100;
#1 $display("%b", po);
# 1  pi=24'b011100010010010001100111;
#1 $display("%b", po);
# 1  pi=24'b111011011101010111111100;
#1 $display("%b", po);
# 1  pi=24'b011111101100101111011101;
#1 $display("%b", po);
# 1  pi=24'b011011010001011101111101;
#1 $display("%b", po);
# 1  pi=24'b001011010001011011101011;
#1 $display("%b", po);
# 1  pi=24'b110100101110011010110010;
#1 $display("%b", po);
# 1  pi=24'b110001111111101100110010;
#1 $display("%b", po);
# 1  pi=24'b011000101100010001100110;
#1 $display("%b", po);
# 1  pi=24'b110011110110111011111010;
#1 $display("%b", po);
# 1  pi=24'b001110101111010010111000;
#1 $display("%b", po);
# 1  pi=24'b100110000101010100110101;
#1 $display("%b", po);
# 1  pi=24'b101111001001011011101110;
#1 $display("%b", po);
# 1  pi=24'b110010011000111010000110;
#1 $display("%b", po);
# 1  pi=24'b000100101000010100011000;
#1 $display("%b", po);
# 1  pi=24'b111100010111111010000101;
#1 $display("%b", po);
# 1  pi=24'b001110101000010010110000;
#1 $display("%b", po);
# 1  pi=24'b100000001000101011010000;
#1 $display("%b", po);
# 1  pi=24'b101001011010111110010010;
#1 $display("%b", po);
# 1  pi=24'b001100000010110010001011;
#1 $display("%b", po);
# 1  pi=24'b110011101011000101100011;
#1 $display("%b", po);
# 1  pi=24'b101110010101010111110001;
#1 $display("%b", po);
# 1  pi=24'b001011100110000110011110;
#1 $display("%b", po);
# 1  pi=24'b110100100101011100101100;
#1 $display("%b", po);
# 1  pi=24'b001000110011011111000011;
#1 $display("%b", po);
# 1  pi=24'b100110000000001000110100;
#1 $display("%b", po);
# 1  pi=24'b001000101111010010001001;
#1 $display("%b", po);
# 1  pi=24'b101001111001100011001110;
#1 $display("%b", po);
# 1  pi=24'b010110101100101110101111;
#1 $display("%b", po);
# 1  pi=24'b111111101101001011100001;
#1 $display("%b", po);
# 1  pi=24'b100101010000100101000101;
#1 $display("%b", po);
# 1  pi=24'b100010101000110100001101;
#1 $display("%b", po);
# 1  pi=24'b010111011110110000101001;
#1 $display("%b", po);
# 1  pi=24'b010101010011101001010000;
#1 $display("%b", po);
# 1  pi=24'b010111100001110000100101;
#1 $display("%b", po);
# 1  pi=24'b100010001100000001000110;
#1 $display("%b", po);
# 1  pi=24'b000011010011010111110000;
#1 $display("%b", po);
# 1  pi=24'b000000110001001010111100;
#1 $display("%b", po);
# 1  pi=24'b111001101010101100100001;
#1 $display("%b", po);
# 1  pi=24'b000111100101011101110011;
#1 $display("%b", po);
# 1  pi=24'b001110110110100000110010;
#1 $display("%b", po);
# 1  pi=24'b111011100100100110111011;
#1 $display("%b", po);
# 1  pi=24'b110001110111101110100010;
#1 $display("%b", po);
# 1  pi=24'b101110110011010000010111;
#1 $display("%b", po);
# 1  pi=24'b001010010000110100110110;
#1 $display("%b", po);
# 1  pi=24'b110000000111000100011001;
#1 $display("%b", po);
# 1  pi=24'b110000000101101000110001;
#1 $display("%b", po);
# 1  pi=24'b101001101101001000011011;
#1 $display("%b", po);
# 1  pi=24'b101000001100000001100100;
#1 $display("%b", po);
# 1  pi=24'b101010001010101100101000;
#1 $display("%b", po);
# 1  pi=24'b011000101111001101111011;
#1 $display("%b", po);
# 1  pi=24'b000011001010010011001000;
#1 $display("%b", po);
# 1  pi=24'b111101110011111110011110;
#1 $display("%b", po);
# 1  pi=24'b111001101110101110110111;
#1 $display("%b", po);
# 1  pi=24'b010101100010101001000011;
#1 $display("%b", po);
# 1  pi=24'b001001000111110010110100;
#1 $display("%b", po);
# 1  pi=24'b010000110010101101111101;
#1 $display("%b", po);
# 1  pi=24'b100011001011011011000011;
#1 $display("%b", po);
# 1  pi=24'b000111010011101000011011;
#1 $display("%b", po);
# 1  pi=24'b111110001011001101100011;
#1 $display("%b", po);
# 1  pi=24'b110111111011100100100000;
#1 $display("%b", po);
# 1  pi=24'b101010100010101001001110;
#1 $display("%b", po);
# 1  pi=24'b001000010111001100000010;
#1 $display("%b", po);
# 1  pi=24'b011111011001000100010110;
#1 $display("%b", po);
# 1  pi=24'b010011001011011000001011;
#1 $display("%b", po);
# 1  pi=24'b111111100111000001010010;
#1 $display("%b", po);
# 1  pi=24'b101100101001010111010111;
#1 $display("%b", po);
# 1  pi=24'b001110001000010100101011;
#1 $display("%b", po);
# 1  pi=24'b110001100100010001100111;
#1 $display("%b", po);
# 1  pi=24'b000111100110100001000000;
#1 $display("%b", po);
# 1  pi=24'b001010000010111101100110;
#1 $display("%b", po);
# 1  pi=24'b111000010111101000000110;
#1 $display("%b", po);
# 1  pi=24'b001010011110001111011010;
#1 $display("%b", po);
# 1  pi=24'b100100011101000110101010;
#1 $display("%b", po);
# 1  pi=24'b101001101101000011000000;
#1 $display("%b", po);
# 1  pi=24'b100101010001101001000110;
#1 $display("%b", po);
# 1  pi=24'b111010000110000110000101;
#1 $display("%b", po);
# 1  pi=24'b010111001001100111100001;
#1 $display("%b", po);
# 1  pi=24'b110111011100000100100001;
#1 $display("%b", po);
# 1  pi=24'b011011101110001001110110;
#1 $display("%b", po);
# 1  pi=24'b010100100101110000011011;
#1 $display("%b", po);
# 1  pi=24'b010000011110001111100010;
#1 $display("%b", po);
# 1  pi=24'b110001001010000000011101;
#1 $display("%b", po);
# 1  pi=24'b111111101000000111100111;
#1 $display("%b", po);
# 1  pi=24'b000100000010010111101101;
#1 $display("%b", po);
# 1  pi=24'b010001101010010011011101;
#1 $display("%b", po);
# 1  pi=24'b101001010110000011001110;
#1 $display("%b", po);
# 1  pi=24'b100000010111110101010000;
#1 $display("%b", po);
# 1  pi=24'b111010011101111001110011;
#1 $display("%b", po);
# 1  pi=24'b001010011001101110011111;
#1 $display("%b", po);
# 1  pi=24'b010010111100011011011011;
#1 $display("%b", po);
# 1  pi=24'b110111111001101100101101;
#1 $display("%b", po);
# 1  pi=24'b000010011001011100100001;
#1 $display("%b", po);
# 1  pi=24'b100011111011010010001011;
#1 $display("%b", po);
# 1  pi=24'b000010101011000011100101;
#1 $display("%b", po);
# 1  pi=24'b001011101010100111010001;
#1 $display("%b", po);
# 1  pi=24'b101010101101110101001111;
#1 $display("%b", po);
# 1  pi=24'b111110111111110000011010;
#1 $display("%b", po);
# 1  pi=24'b010111110101010100110010;
#1 $display("%b", po);
# 1  pi=24'b010000110111011001100010;
#1 $display("%b", po);
# 1  pi=24'b111110001010101010000101;
#1 $display("%b", po);
# 1  pi=24'b011011001111000000000111;
#1 $display("%b", po);
# 1  pi=24'b100011111011111101110110;
#1 $display("%b", po);
# 1  pi=24'b001010011000110000110100;
#1 $display("%b", po);
# 1  pi=24'b011011111110101011001000;
#1 $display("%b", po);
# 1  pi=24'b011100111101011000100010;
#1 $display("%b", po);
# 1  pi=24'b010100001101000010111010;
#1 $display("%b", po);
# 1  pi=24'b000101111101010010111111;
#1 $display("%b", po);
# 1  pi=24'b010111110110000000100100;
#1 $display("%b", po);
# 1  pi=24'b000010101011011001000100;
#1 $display("%b", po);
# 1  pi=24'b101001001110110110110010;
#1 $display("%b", po);
# 1  pi=24'b011001000101111100110101;
#1 $display("%b", po);
# 1  pi=24'b010010011010000000000111;
#1 $display("%b", po);
# 1  pi=24'b110111101100100001100111;
#1 $display("%b", po);
# 1  pi=24'b010011000000111101001000;
#1 $display("%b", po);
# 1  pi=24'b000001001011000100010011;
#1 $display("%b", po);
# 1  pi=24'b000011110110100111010000;
#1 $display("%b", po);
# 1  pi=24'b010101001011110110101111;
#1 $display("%b", po);
# 1  pi=24'b110101111111011000101111;
#1 $display("%b", po);
# 1  pi=24'b011011110001011001111100;
#1 $display("%b", po);
# 1  pi=24'b110110100110010101100101;
#1 $display("%b", po);
# 1  pi=24'b110011001101010101011111;
#1 $display("%b", po);
# 1  pi=24'b010101101001011101011101;
#1 $display("%b", po);
# 1  pi=24'b000011000101010110101001;
#1 $display("%b", po);
# 1  pi=24'b111000011011110000110010;
#1 $display("%b", po);
# 1  pi=24'b001110111111001000111110;
#1 $display("%b", po);
# 1  pi=24'b111000100001011011011000;
#1 $display("%b", po);
# 1  pi=24'b101011001011100100100010;
#1 $display("%b", po);
# 1  pi=24'b100011111011101100011110;
#1 $display("%b", po);
# 1  pi=24'b100000101000101011010101;
#1 $display("%b", po);
# 1  pi=24'b001110101100000001010101;
#1 $display("%b", po);
# 1  pi=24'b101011001100110111010111;
#1 $display("%b", po);
# 1  pi=24'b101101011011000100000100;
#1 $display("%b", po);
# 1  pi=24'b110100110111111010011001;
#1 $display("%b", po);
# 1  pi=24'b000111110101100001000110;
#1 $display("%b", po);
# 1  pi=24'b000101111111000110101100;
#1 $display("%b", po);
# 1  pi=24'b101110110110101111011010;
#1 $display("%b", po);
# 1  pi=24'b111011100100001001001100;
#1 $display("%b", po);
# 1  pi=24'b100101111000100111110111;
#1 $display("%b", po);
# 1  pi=24'b001110000100101011111011;
#1 $display("%b", po);
# 1  pi=24'b100101010110110001100011;
#1 $display("%b", po);
# 1  pi=24'b100010111110001111011001;
#1 $display("%b", po);
# 1  pi=24'b010110100100000011101111;
#1 $display("%b", po);
# 1  pi=24'b011001000110000010000010;
#1 $display("%b", po);
# 1  pi=24'b100110101000000100010111;
#1 $display("%b", po);
# 1  pi=24'b100000101010100100010110;
#1 $display("%b", po);
# 1  pi=24'b011110011000110010100000;
#1 $display("%b", po);
# 1  pi=24'b000010100001001101011111;
#1 $display("%b", po);
# 1  pi=24'b100101100101100101101100;
#1 $display("%b", po);
# 1  pi=24'b000101000011101101111111;
#1 $display("%b", po);
# 1  pi=24'b001111001010110100111000;
#1 $display("%b", po);
# 1  pi=24'b011001111110011010010011;
#1 $display("%b", po);
# 1  pi=24'b110110110100011110111010;
#1 $display("%b", po);
# 1  pi=24'b111011011110001011100000;
#1 $display("%b", po);
# 1  pi=24'b001010000101100100100000;
#1 $display("%b", po);
# 1  pi=24'b110101101111110101111111;
#1 $display("%b", po);
# 1  pi=24'b010000010111000001101010;
#1 $display("%b", po);
# 1  pi=24'b011100111100110110000101;
#1 $display("%b", po);
# 1  pi=24'b101111010111011001100101;
#1 $display("%b", po);
# 1  pi=24'b011110011111101100000101;
#1 $display("%b", po);
# 1  pi=24'b110110101001010101111010;
#1 $display("%b", po);
# 1  pi=24'b110011110101110110110001;
#1 $display("%b", po);
# 1  pi=24'b100100010001000110111011;
#1 $display("%b", po);
# 1  pi=24'b101011100001100100111010;
#1 $display("%b", po);
# 1  pi=24'b001001111000110010000011;
#1 $display("%b", po);
# 1  pi=24'b111110100001101000000011;
#1 $display("%b", po);
# 1  pi=24'b100010011010011110011010;
#1 $display("%b", po);
# 1  pi=24'b000111001110101100010111;
#1 $display("%b", po);
# 1  pi=24'b111110100111011011000111;
#1 $display("%b", po);
# 1  pi=24'b001010011111101001010100;
#1 $display("%b", po);
# 1  pi=24'b001001110110100111101011;
#1 $display("%b", po);
# 1  pi=24'b101000110110100001001111;
#1 $display("%b", po);
# 1  pi=24'b001100010100001100101101;
#1 $display("%b", po);
# 1  pi=24'b110000011000101010001100;
#1 $display("%b", po);
# 1  pi=24'b100111011111101110001000;
#1 $display("%b", po);
# 1  pi=24'b101000100111111011101000;
#1 $display("%b", po);
# 1  pi=24'b100100010000011011111111;
#1 $display("%b", po);
# 1  pi=24'b010101111111110000110010;
#1 $display("%b", po);
# 1  pi=24'b111110101011100111110001;
#1 $display("%b", po);
# 1  pi=24'b001010111100101000101000;
#1 $display("%b", po);
# 1  pi=24'b011110000110010010101100;
#1 $display("%b", po);
# 1  pi=24'b110111000110100011000010;
#1 $display("%b", po);
# 1  pi=24'b100000001101110111111010;
#1 $display("%b", po);
# 1  pi=24'b011011000000000001011101;
#1 $display("%b", po);
# 1  pi=24'b110011111101011111011100;
#1 $display("%b", po);
# 1  pi=24'b001010001010011111101110;
#1 $display("%b", po);
# 1  pi=24'b010111010110110011111111;
#1 $display("%b", po);
# 1  pi=24'b111000101000010001100100;
#1 $display("%b", po);
# 1  pi=24'b100001111010011101111101;
#1 $display("%b", po);
# 1  pi=24'b000011011111001010110111;
#1 $display("%b", po);
# 1  pi=24'b110001110110010011011010;
#1 $display("%b", po);
# 1  pi=24'b011001110010101001001110;
#1 $display("%b", po);
# 1  pi=24'b111001101101100101111001;
#1 $display("%b", po);
# 1  pi=24'b100010001110100110010000;
#1 $display("%b", po);
# 1  pi=24'b011101101111000111000000;
#1 $display("%b", po);
# 1  pi=24'b100100100111010010010111;
#1 $display("%b", po);
# 1  pi=24'b010000000000001010011111;
#1 $display("%b", po);
# 1  pi=24'b010111010101111100011100;
#1 $display("%b", po);
# 1  pi=24'b010010101110101111010101;
#1 $display("%b", po);
# 1  pi=24'b000010010101011001001010;
#1 $display("%b", po);
# 1  pi=24'b001001101101111011110000;
#1 $display("%b", po);
# 1  pi=24'b000101000101111011100010;
#1 $display("%b", po);
# 1  pi=24'b011101100110010110011111;
#1 $display("%b", po);
# 1  pi=24'b101111010010101101010100;
#1 $display("%b", po);
# 1  pi=24'b110011001000111101000011;
#1 $display("%b", po);
# 1  pi=24'b101110000111111101100010;
#1 $display("%b", po);
# 1  pi=24'b011001111110101110001000;
#1 $display("%b", po);
# 1  pi=24'b110001111010100001001101;
#1 $display("%b", po);
# 1  pi=24'b001100100111110000110011;
#1 $display("%b", po);
# 1  pi=24'b011110100111000011001110;
#1 $display("%b", po);
# 1  pi=24'b001101000100110000001001;
#1 $display("%b", po);
# 1  pi=24'b011001111110111010000011;
#1 $display("%b", po);
# 1  pi=24'b010100000101001001100110;
#1 $display("%b", po);
# 1  pi=24'b111011011001101101111010;
#1 $display("%b", po);
# 1  pi=24'b111000000101000101100000;
#1 $display("%b", po);
# 1  pi=24'b100100011001111111010100;
#1 $display("%b", po);
# 1  pi=24'b111001110100110100001110;
#1 $display("%b", po);
# 1  pi=24'b001100101100111100000001;
#1 $display("%b", po);
# 1  pi=24'b010000001101000010101000;
#1 $display("%b", po);
# 1  pi=24'b010011110101110010011010;
#1 $display("%b", po);
# 1  pi=24'b111100100100111100001100;
#1 $display("%b", po);
# 1  pi=24'b101011110100010000110111;
#1 $display("%b", po);
# 1  pi=24'b110011110101100111010100;
#1 $display("%b", po);
# 1  pi=24'b111000111111000010001010;
#1 $display("%b", po);
# 1  pi=24'b001110101000100011111111;
#1 $display("%b", po);
# 1  pi=24'b001101101001111000011000;
#1 $display("%b", po);
# 1  pi=24'b101011100010101110001001;
#1 $display("%b", po);
# 1  pi=24'b110010001010011011010111;
#1 $display("%b", po);
# 1  pi=24'b101001111000011011111011;
#1 $display("%b", po);
# 1  pi=24'b100100111111010101001001;
#1 $display("%b", po);
# 1  pi=24'b110100110111000110111110;
#1 $display("%b", po);
# 1  pi=24'b001101100001010100101000;
#1 $display("%b", po);
# 1  pi=24'b110010110100010100001011;
#1 $display("%b", po);
# 1  pi=24'b100110111110101000101010;
#1 $display("%b", po);
# 1  pi=24'b011011110011010110101110;
#1 $display("%b", po);
# 1  pi=24'b001111101010101000100010;
#1 $display("%b", po);
# 1  pi=24'b001101101000110101101100;
#1 $display("%b", po);
# 1  pi=24'b001000010010001101001011;
#1 $display("%b", po);
# 1  pi=24'b100111110111101001111101;
#1 $display("%b", po);
# 1  pi=24'b011001011000101101010000;
#1 $display("%b", po);
# 1  pi=24'b111111111111001101011110;
#1 $display("%b", po);
# 1  pi=24'b111011011110100000110010;
#1 $display("%b", po);
# 1  pi=24'b100111101101100010101001;
#1 $display("%b", po);
# 1  pi=24'b111010001100000000010101;
#1 $display("%b", po);
# 1  pi=24'b101100011111100111101010;
#1 $display("%b", po);
# 1  pi=24'b101001111011010101101010;
#1 $display("%b", po);
# 1  pi=24'b000011100111100110100001;
#1 $display("%b", po);
# 1  pi=24'b101010011001110110111101;
#1 $display("%b", po);
# 1  pi=24'b010110011010110010110101;
#1 $display("%b", po);
# 1  pi=24'b011001101110110011001010;
#1 $display("%b", po);
# 1  pi=24'b011000101000110110001011;
#1 $display("%b", po);
# 1  pi=24'b001111111101110000001101;
#1 $display("%b", po);
# 1  pi=24'b110111101011101001001101;
#1 $display("%b", po);
# 1  pi=24'b110100010001001101001101;
#1 $display("%b", po);
# 1  pi=24'b101010110010111001001000;
#1 $display("%b", po);
# 1  pi=24'b111001010010010011001011;
#1 $display("%b", po);
# 1  pi=24'b000101000011101111110010;
#1 $display("%b", po);
# 1  pi=24'b101000001010110110011000;
#1 $display("%b", po);
# 1  pi=24'b100010110100001010110100;
#1 $display("%b", po);
# 1  pi=24'b011111111000100001011000;
#1 $display("%b", po);
# 1  pi=24'b010110011101110110001001;
#1 $display("%b", po);
# 1  pi=24'b100000100001100111101010;
#1 $display("%b", po);
# 1  pi=24'b101000111110111000111001;
#1 $display("%b", po);
# 1  pi=24'b001000110110011010101100;
#1 $display("%b", po);
# 1  pi=24'b010100000110010011010100;
#1 $display("%b", po);
# 1  pi=24'b110000011110001000111000;
#1 $display("%b", po);
# 1  pi=24'b110111000001011011101010;
#1 $display("%b", po);
# 1  pi=24'b001111101110100000011011;
#1 $display("%b", po);
# 1  pi=24'b100111011001001010110101;
#1 $display("%b", po);
# 1  pi=24'b110101101000110000110100;
#1 $display("%b", po);
# 1  pi=24'b101110010111011011011010;
#1 $display("%b", po);
# 1  pi=24'b111000110001000011000101;
#1 $display("%b", po);
# 1  pi=24'b101110011001100111000111;
#1 $display("%b", po);
# 1  pi=24'b010000010110011111101110;
#1 $display("%b", po);
# 1  pi=24'b110101000110110101100011;
#1 $display("%b", po);
# 1  pi=24'b010110011000110011011110;
#1 $display("%b", po);
# 1  pi=24'b111001110110111101110010;
#1 $display("%b", po);
# 1  pi=24'b101110001011010101011110;
#1 $display("%b", po);
# 1  pi=24'b010110010101110010101101;
#1 $display("%b", po);
# 1  pi=24'b010011101111100010011110;
#1 $display("%b", po);
# 1  pi=24'b101101010111111101011010;
#1 $display("%b", po);
# 1  pi=24'b000010111111000100011110;
#1 $display("%b", po);
# 1  pi=24'b101111111111010100110111;
#1 $display("%b", po);
# 1  pi=24'b011001010001000111001101;
#1 $display("%b", po);
# 1  pi=24'b000011000100101110010100;
#1 $display("%b", po);
# 1  pi=24'b000100010001000110011001;
#1 $display("%b", po);
# 1  pi=24'b110011010101110110111101;
#1 $display("%b", po);
# 1  pi=24'b110000001010111100000110;
#1 $display("%b", po);
# 1  pi=24'b111111100110010011000111;
#1 $display("%b", po);
# 1  pi=24'b111001000111100010101000;
#1 $display("%b", po);
# 1  pi=24'b011010101111010011010001;
#1 $display("%b", po);
# 1  pi=24'b010111010011110011111011;
#1 $display("%b", po);
# 1  pi=24'b101011010000001000010110;
#1 $display("%b", po);
# 1  pi=24'b000101110000001110000101;
#1 $display("%b", po);
# 1  pi=24'b001101101010000110101110;
#1 $display("%b", po);
# 1  pi=24'b010000100111110001010110;
#1 $display("%b", po);
# 1  pi=24'b111011111110000011000011;
#1 $display("%b", po);
# 1  pi=24'b111011100110110100011110;
#1 $display("%b", po);
# 1  pi=24'b001110001000011111101011;
#1 $display("%b", po);
# 1  pi=24'b100111011111001111101011;
#1 $display("%b", po);
# 1  pi=24'b110001101110001000111101;
#1 $display("%b", po);
# 1  pi=24'b001001010111010111101101;
#1 $display("%b", po);
# 1  pi=24'b100110100001001001010111;
#1 $display("%b", po);
# 1  pi=24'b110111100010110111011010;
#1 $display("%b", po);
# 1  pi=24'b101011001011100111000110;
#1 $display("%b", po);
# 1  pi=24'b000000110100001100101111;
#1 $display("%b", po);
# 1  pi=24'b001110111111111110110011;
#1 $display("%b", po);
# 1  pi=24'b011001000101010110100111;
#1 $display("%b", po);
# 1  pi=24'b111100001011111101001100;
#1 $display("%b", po);
# 1  pi=24'b010111110100110011110101;
#1 $display("%b", po);
# 1  pi=24'b100101000110100011000010;
#1 $display("%b", po);
# 1  pi=24'b101110010101101010101011;
#1 $display("%b", po);
# 1  pi=24'b101011101100000101011011;
#1 $display("%b", po);
# 1  pi=24'b001000100001110111000000;
#1 $display("%b", po);
# 1  pi=24'b001010001001100100011000;
#1 $display("%b", po);
# 1  pi=24'b000101100010101110111010;
#1 $display("%b", po);
# 1  pi=24'b001001111000011001011011;
#1 $display("%b", po);
# 1  pi=24'b100111100111100100110011;
#1 $display("%b", po);
# 1  pi=24'b110101000110010001100111;
#1 $display("%b", po);
# 1  pi=24'b000001100110110011111010;
#1 $display("%b", po);
# 1  pi=24'b010101101101101001101011;
#1 $display("%b", po);
# 1  pi=24'b011110010000111110100111;
#1 $display("%b", po);
# 1  pi=24'b101011110011101110110000;
#1 $display("%b", po);
# 1  pi=24'b000101010011111101000011;
#1 $display("%b", po);
# 1  pi=24'b101101001011110100011100;
#1 $display("%b", po);
# 1  pi=24'b111000001000101111101111;
#1 $display("%b", po);
# 1  pi=24'b010100101011110100001010;
#1 $display("%b", po);
# 1  pi=24'b101111110101100111100100;
#1 $display("%b", po);
# 1  pi=24'b000011001110000001010001;
#1 $display("%b", po);
# 1  pi=24'b011000110000111011110011;
#1 $display("%b", po);
# 1  pi=24'b101111001110001111010100;
#1 $display("%b", po);
# 1  pi=24'b010000111110111110000001;
#1 $display("%b", po);
# 1  pi=24'b000010000000101101101110;
#1 $display("%b", po);
# 1  pi=24'b010000101001100010101111;
#1 $display("%b", po);
# 1  pi=24'b110001000010000110011101;
#1 $display("%b", po);
# 1  pi=24'b111011001101100101011011;
#1 $display("%b", po);
# 1  pi=24'b101100000000010101101101;
#1 $display("%b", po);
# 1  pi=24'b101101011101001011101000;
#1 $display("%b", po);
# 1  pi=24'b110011001110111110101111;
#1 $display("%b", po);
# 1  pi=24'b111111010101000111011100;
#1 $display("%b", po);
# 1  pi=24'b011001110101100011001001;
#1 $display("%b", po);
# 1  pi=24'b010001110111110011010111;
#1 $display("%b", po);
# 1  pi=24'b111011111001100001100010;
#1 $display("%b", po);
# 1  pi=24'b100101101111011000000010;
#1 $display("%b", po);
# 1  pi=24'b000110110111011111110000;
#1 $display("%b", po);
# 1  pi=24'b000110111000100111100001;
#1 $display("%b", po);
# 1  pi=24'b110111011001011111000000;
#1 $display("%b", po);
# 1  pi=24'b011000100000010001000110;
#1 $display("%b", po);
# 1  pi=24'b010111010111011011100011;
#1 $display("%b", po);
# 1  pi=24'b011100010111000010010110;
#1 $display("%b", po);
# 1  pi=24'b111011011100000110001001;
#1 $display("%b", po);
# 1  pi=24'b111010000110101101001010;
#1 $display("%b", po);
# 1  pi=24'b011000100101101101011010;
#1 $display("%b", po);
# 1  pi=24'b100000011100000011011011;
#1 $display("%b", po);
# 1  pi=24'b000010011001011000010100;
#1 $display("%b", po);
# 1  pi=24'b110000101001000100100010;
#1 $display("%b", po);
# 1  pi=24'b010011101111001100111110;
#1 $display("%b", po);
# 1  pi=24'b101100000010110101111100;
#1 $display("%b", po);
# 1  pi=24'b001010101011100000011111;
#1 $display("%b", po);
# 1  pi=24'b100010000001101011000010;
#1 $display("%b", po);
# 1  pi=24'b000111001100001000001010;
#1 $display("%b", po);
# 1  pi=24'b000001111000000001110011;
#1 $display("%b", po);
# 1  pi=24'b111001011100001001001000;
#1 $display("%b", po);
# 1  pi=24'b010001111111001010110100;
#1 $display("%b", po);
# 1  pi=24'b011111110001010011001101;
#1 $display("%b", po);
# 1  pi=24'b100100111010000101000101;
#1 $display("%b", po);
# 1  pi=24'b100001000110101011110110;
#1 $display("%b", po);
# 1  pi=24'b110110100100001011101101;
#1 $display("%b", po);
# 1  pi=24'b110011111100100001101101;
#1 $display("%b", po);
# 1  pi=24'b111010111101000100111010;
#1 $display("%b", po);
# 1  pi=24'b000111000101101100100001;
#1 $display("%b", po);
# 1  pi=24'b100011101001001111111111;
#1 $display("%b", po);
# 1  pi=24'b111100110010111101111101;
#1 $display("%b", po);
# 1  pi=24'b010010111000101110001001;
#1 $display("%b", po);
# 1  pi=24'b111111001000011000001000;
#1 $display("%b", po);
# 1  pi=24'b101001111100100000111011;
#1 $display("%b", po);
# 1  pi=24'b000101000001011110011011;
#1 $display("%b", po);
# 1  pi=24'b111001101101111010101111;
#1 $display("%b", po);
# 1  pi=24'b010000100000100110100111;
#1 $display("%b", po);
# 1  pi=24'b101010100101010110110101;
#1 $display("%b", po);
# 1  pi=24'b000110111100111011011110;
#1 $display("%b", po);
# 1  pi=24'b010001011000000100000100;
#1 $display("%b", po);
# 1  pi=24'b111010010010111111100100;
#1 $display("%b", po);
# 1  pi=24'b100110010001011110010000;
#1 $display("%b", po);
# 1  pi=24'b011111001111101111001111;
#1 $display("%b", po);
# 1  pi=24'b010101110011110101000000;
#1 $display("%b", po);
# 1  pi=24'b100101101000100010001001;
#1 $display("%b", po);
# 1  pi=24'b010100001101001110100101;
#1 $display("%b", po);
# 1  pi=24'b001100111000011011000001;
#1 $display("%b", po);
# 1  pi=24'b011110110001000101000101;
#1 $display("%b", po);
# 1  pi=24'b111000010100111110000001;
#1 $display("%b", po);
# 1  pi=24'b110101101011100101001111;
#1 $display("%b", po);
# 1  pi=24'b100110101101110001111101;
#1 $display("%b", po);
# 1  pi=24'b111000010110110001101111;
#1 $display("%b", po);
# 1  pi=24'b111110110001001000011010;
#1 $display("%b", po);
# 1  pi=24'b001010001011011001011010;
#1 $display("%b", po);
# 1  pi=24'b110010010111010001000101;
#1 $display("%b", po);
# 1  pi=24'b000100011100001011110110;
#1 $display("%b", po);
# 1  pi=24'b011011000110010110111000;
#1 $display("%b", po);
# 1  pi=24'b011110110101001001100001;
#1 $display("%b", po);
# 1  pi=24'b101000010001101001110010;
#1 $display("%b", po);
# 1  pi=24'b101110000010011110001100;
#1 $display("%b", po);
# 1  pi=24'b110011010011011000110000;
#1 $display("%b", po);
# 1  pi=24'b001011001111111010101001;
#1 $display("%b", po);
# 1  pi=24'b111100111100010101011010;
#1 $display("%b", po);
# 1  pi=24'b001110110100001001100001;
#1 $display("%b", po);
# 1  pi=24'b111010100011110000011111;
#1 $display("%b", po);
# 1  pi=24'b010101001110011101111101;
#1 $display("%b", po);
# 1  pi=24'b100101101000110000011100;
#1 $display("%b", po);
# 1  pi=24'b100110011000100111000011;
#1 $display("%b", po);
# 1  pi=24'b000000101111001110111110;
#1 $display("%b", po);
# 1  pi=24'b111011011100000010000010;
#1 $display("%b", po);
# 1  pi=24'b001101100011011011000001;
#1 $display("%b", po);
# 1  pi=24'b111110100010100000111111;
#1 $display("%b", po);
# 1  pi=24'b000100011100001010101100;
#1 $display("%b", po);
# 1  pi=24'b110110111101010000100000;
#1 $display("%b", po);
# 1  pi=24'b000010111100001101011000;
#1 $display("%b", po);
# 1  pi=24'b011100111000110101100000;
#1 $display("%b", po);
# 1  pi=24'b100010000111011110010111;
#1 $display("%b", po);
# 1  pi=24'b011010010000100001111101;
#1 $display("%b", po);
# 1  pi=24'b010101101011111001111011;
#1 $display("%b", po);
# 1  pi=24'b001111111101110001000010;
#1 $display("%b", po);
# 1  pi=24'b111011010101100111110001;
#1 $display("%b", po);
# 1  pi=24'b111110001111100101001101;
#1 $display("%b", po);
# 1  pi=24'b000111111011111001010000;
#1 $display("%b", po);
# 1  pi=24'b010001110111100001100110;
#1 $display("%b", po);
# 1  pi=24'b000001000101100110001101;
#1 $display("%b", po);
# 1  pi=24'b000000101110001100000001;
#1 $display("%b", po);
# 1  pi=24'b110000111111011000110110;
#1 $display("%b", po);
# 1  pi=24'b101111101111101011110001;
#1 $display("%b", po);
# 1  pi=24'b010110001110110111000100;
#1 $display("%b", po);
# 1  pi=24'b100111101000010010101111;
#1 $display("%b", po);
# 1  pi=24'b000010001110111100001001;
#1 $display("%b", po);
# 1  pi=24'b001010100101100011000101;
#1 $display("%b", po);
# 1  pi=24'b101001000001101110011001;
#1 $display("%b", po);
# 1  pi=24'b011011100011001101111110;
#1 $display("%b", po);
# 1  pi=24'b000101111110100101111110;
#1 $display("%b", po);
# 1  pi=24'b010011100000100110101101;
#1 $display("%b", po);
# 1  pi=24'b101101001011000101100000;
#1 $display("%b", po);
# 1  pi=24'b010000000010101100100000;
#1 $display("%b", po);
# 1  pi=24'b111110010000100010100010;
#1 $display("%b", po);
# 1  pi=24'b000100010110011111000000;
#1 $display("%b", po);
# 1  pi=24'b010100010001101101000111;
#1 $display("%b", po);
# 1  pi=24'b100010010001011011011011;
#1 $display("%b", po);
# 1  pi=24'b110001001100110111110001;
#1 $display("%b", po);
# 1  pi=24'b010100111000100110100110;
#1 $display("%b", po);
# 1  pi=24'b011110110101000101111100;
#1 $display("%b", po);
# 1  pi=24'b000001010111100111011110;
#1 $display("%b", po);
# 1  pi=24'b111100011011001100100111;
#1 $display("%b", po);
# 1  pi=24'b000100101111100100001010;
#1 $display("%b", po);
# 1  pi=24'b011111010100110011100011;
#1 $display("%b", po);
# 1  pi=24'b110111101010000111101011;
#1 $display("%b", po);
# 1  pi=24'b100000111000101000000111;
#1 $display("%b", po);
# 1  pi=24'b011101100011000000011111;
#1 $display("%b", po);
# 1  pi=24'b011100101100010111110100;
#1 $display("%b", po);
# 1  pi=24'b110000100010101000011111;
#1 $display("%b", po);
# 1  pi=24'b110001110000101110111001;
#1 $display("%b", po);
# 1  pi=24'b011110011000110011011011;
#1 $display("%b", po);
# 1  pi=24'b111111110001000101011111;
#1 $display("%b", po);
# 1  pi=24'b100011000000101010001110;
#1 $display("%b", po);
# 1  pi=24'b010101000000101100111000;
#1 $display("%b", po);
# 1  pi=24'b000111110000101010010000;
#1 $display("%b", po);
# 1  pi=24'b101111000101101100001011;
#1 $display("%b", po);
# 1  pi=24'b001000000001001011110000;
#1 $display("%b", po);
# 1  pi=24'b001111001100000110011010;
#1 $display("%b", po);
# 1  pi=24'b010000001010100100100101;
#1 $display("%b", po);
# 1  pi=24'b011100111010001101000110;
#1 $display("%b", po);
# 1  pi=24'b010111111011100011001110;
#1 $display("%b", po);
# 1  pi=24'b101111110101100100110000;
#1 $display("%b", po);
# 1  pi=24'b110010010011010100001110;
#1 $display("%b", po);
# 1  pi=24'b010111010000000110101101;
#1 $display("%b", po);
# 1  pi=24'b100100110101001010100111;
#1 $display("%b", po);
# 1  pi=24'b110110001101110011111101;
#1 $display("%b", po);
# 1  pi=24'b010100010011111101100000;
#1 $display("%b", po);
# 1  pi=24'b111011111110010110011011;
#1 $display("%b", po);
# 1  pi=24'b101011100001100101011101;
#1 $display("%b", po);
# 1  pi=24'b110010100010101011111000;
#1 $display("%b", po);
# 1  pi=24'b101010100111011110010111;
#1 $display("%b", po);
# 1  pi=24'b101011100010011111000101;
#1 $display("%b", po);
# 1  pi=24'b011001100111101011111110;
#1 $display("%b", po);
# 1  pi=24'b101101101111110110011110;
#1 $display("%b", po);
# 1  pi=24'b001010001011011000000111;
#1 $display("%b", po);
# 1  pi=24'b001010011111110010101100;
#1 $display("%b", po);
# 1  pi=24'b110000101010110001000111;
#1 $display("%b", po);
# 1  pi=24'b010101111110111111011011;
#1 $display("%b", po);
# 1  pi=24'b100101011101101000100000;
#1 $display("%b", po);
# 1  pi=24'b101100001000010111111001;
#1 $display("%b", po);
# 1  pi=24'b001010111000000001111000;
#1 $display("%b", po);
# 1  pi=24'b001001100111011000101110;
#1 $display("%b", po);
# 1  pi=24'b100000011010101011001111;
#1 $display("%b", po);
# 1  pi=24'b111011101100100111000001;
#1 $display("%b", po);
# 1  pi=24'b111001101011011111101111;
#1 $display("%b", po);
# 1  pi=24'b011100011110110101001010;
#1 $display("%b", po);
# 1  pi=24'b101011011101100101010000;
#1 $display("%b", po);
# 1  pi=24'b110001100110001100001001;
#1 $display("%b", po);
# 1  pi=24'b111111000010011101100111;
#1 $display("%b", po);
# 1  pi=24'b111010101000010111101000;
#1 $display("%b", po);
# 1  pi=24'b011001010001011101000101;
#1 $display("%b", po);
# 1  pi=24'b010010100010000000000011;
#1 $display("%b", po);
# 1  pi=24'b110101101000010001010010;
#1 $display("%b", po);
# 1  pi=24'b110001101111110000101111;
#1 $display("%b", po);
# 1  pi=24'b001001110101000110000101;
#1 $display("%b", po);
# 1  pi=24'b000111010011001111001010;
#1 $display("%b", po);
# 1  pi=24'b000010101101110010010001;
#1 $display("%b", po);
# 1  pi=24'b101001100010110001001100;
#1 $display("%b", po);
# 1  pi=24'b100010011100100000000110;
#1 $display("%b", po);
# 1  pi=24'b110111110011000000111111;
#1 $display("%b", po);
# 1  pi=24'b001001001111100101111101;
#1 $display("%b", po);
# 1  pi=24'b000111100111000000111111;
#1 $display("%b", po);
# 1  pi=24'b110010001110001000100111;
#1 $display("%b", po);
# 1  pi=24'b001101100000101100110000;
#1 $display("%b", po);
# 1  pi=24'b100101011011100010010001;
#1 $display("%b", po);
# 1  pi=24'b010011100000110110000000;
#1 $display("%b", po);
# 1  pi=24'b000001100000101011100011;
#1 $display("%b", po);
# 1  pi=24'b101011011001101001001000;
#1 $display("%b", po);
# 1  pi=24'b100000010001111110000101;
#1 $display("%b", po);
# 1  pi=24'b111110101100100001001110;
#1 $display("%b", po);
# 1  pi=24'b000100011110100000010101;
#1 $display("%b", po);
# 1  pi=24'b010001011100111111010100;
#1 $display("%b", po);
# 1  pi=24'b101001110011011101001011;
#1 $display("%b", po);
# 1  pi=24'b100011000000101100100110;
#1 $display("%b", po);
# 1  pi=24'b010011001101011001100011;
#1 $display("%b", po);
# 1  pi=24'b101000001001010000100011;
#1 $display("%b", po);
# 1  pi=24'b011111111100110101000101;
#1 $display("%b", po);
# 1  pi=24'b000010010100000110111100;
#1 $display("%b", po);
# 1  pi=24'b000010111101001111011011;
#1 $display("%b", po);
# 1  pi=24'b100000011011100110110010;
#1 $display("%b", po);
# 1  pi=24'b100110110100010111000011;
#1 $display("%b", po);
# 1  pi=24'b011101101010011101110000;
#1 $display("%b", po);
# 1  pi=24'b010101000011011001100100;
#1 $display("%b", po);
# 1  pi=24'b111100100001110011111011;
#1 $display("%b", po);
# 1  pi=24'b001001101101110001010000;
#1 $display("%b", po);
# 1  pi=24'b000010111011001101011001;
#1 $display("%b", po);
# 1  pi=24'b110100101111000010100100;
#1 $display("%b", po);
# 1  pi=24'b101010000010101001010011;
#1 $display("%b", po);
# 1  pi=24'b100111010001100011011010;
#1 $display("%b", po);
# 1  pi=24'b101011110011010100101010;
#1 $display("%b", po);
# 1  pi=24'b100111010000100001000101;
#1 $display("%b", po);
# 1  pi=24'b011000011100001110101011;
#1 $display("%b", po);
# 1  pi=24'b001011011111000101101111;
#1 $display("%b", po);
# 1  pi=24'b001001110001001100011000;
#1 $display("%b", po);
# 1  pi=24'b010000011011011111010001;
#1 $display("%b", po);
# 1  pi=24'b011010111010101110010111;
#1 $display("%b", po);
# 1  pi=24'b111111101010101100011010;
#1 $display("%b", po);
# 1  pi=24'b101011111111000111101011;
#1 $display("%b", po);
# 1  pi=24'b101100101101010111011010;
#1 $display("%b", po);
# 1  pi=24'b110000001110100100011100;
#1 $display("%b", po);
# 1  pi=24'b000110100111011010001101;
#1 $display("%b", po);
# 1  pi=24'b010101010010011001000111;
#1 $display("%b", po);
# 1  pi=24'b101100111101011111100011;
#1 $display("%b", po);
# 1  pi=24'b010001111111000110101010;
#1 $display("%b", po);
# 1  pi=24'b101110111110100101111111;
#1 $display("%b", po);
# 1  pi=24'b100001000011110011110100;
#1 $display("%b", po);
# 1  pi=24'b011110100001001001011101;
#1 $display("%b", po);
# 1  pi=24'b101111010011101000001000;
#1 $display("%b", po);
# 1  pi=24'b101100010101110001100100;
#1 $display("%b", po);
# 1  pi=24'b110011111000001100001000;
#1 $display("%b", po);
# 1  pi=24'b100011000100010001111100;
#1 $display("%b", po);
# 1  pi=24'b100011110101000011111000;
#1 $display("%b", po);
# 1  pi=24'b101110100100010000001111;
#1 $display("%b", po);
# 1  pi=24'b101110111001100100100111;
#1 $display("%b", po);
# 1  pi=24'b010000000110011000000101;
#1 $display("%b", po);
# 1  pi=24'b001011110011110101000101;
#1 $display("%b", po);
# 1  pi=24'b101100001000010000101100;
#1 $display("%b", po);
# 1  pi=24'b111100000111011101110101;
#1 $display("%b", po);
# 1  pi=24'b100110110011101101011000;
#1 $display("%b", po);
# 1  pi=24'b010100101101011000010010;
#1 $display("%b", po);
# 1  pi=24'b111001000100001000101000;
#1 $display("%b", po);
# 1  pi=24'b000100100110100010000010;
#1 $display("%b", po);
# 1  pi=24'b100101010110101100100000;
#1 $display("%b", po);
# 1  pi=24'b100011011111000011111101;
#1 $display("%b", po);
# 1  pi=24'b001101100111011110000100;
#1 $display("%b", po);
# 1  pi=24'b000011110111000111010000;
#1 $display("%b", po);
# 1  pi=24'b110010110000001111011001;
#1 $display("%b", po);
# 1  pi=24'b010110111011100011000101;
#1 $display("%b", po);
# 1  pi=24'b110011101111101101111011;
#1 $display("%b", po);
# 1  pi=24'b000011011110101010000100;
#1 $display("%b", po);
# 1  pi=24'b011110010111100011100011;
#1 $display("%b", po);
# 1  pi=24'b000111011111011000111101;
#1 $display("%b", po);
# 1  pi=24'b011100110111100110001010;
#1 $display("%b", po);
# 1  pi=24'b100110000111100101110110;
#1 $display("%b", po);
# 1  pi=24'b110110111010001101010011;
#1 $display("%b", po);
# 1  pi=24'b110010100001010101011101;
#1 $display("%b", po);
# 1  pi=24'b000011011011011010110100;
#1 $display("%b", po);
# 1  pi=24'b010110111000001110000011;
#1 $display("%b", po);
# 1  pi=24'b010101110100001010100110;
#1 $display("%b", po);
# 1  pi=24'b100010110101000011111110;
#1 $display("%b", po);
# 1  pi=24'b100000110101010000101100;
#1 $display("%b", po);
# 1  pi=24'b101111101000000100100111;
#1 $display("%b", po);
# 1  pi=24'b100001100111100011100110;
#1 $display("%b", po);
# 1  pi=24'b110111011110110111111100;
#1 $display("%b", po);
# 1  pi=24'b011001010111000101111010;
#1 $display("%b", po);
# 1  pi=24'b101010011101010000010100;
#1 $display("%b", po);
# 1  pi=24'b111001110001001101001001;
#1 $display("%b", po);
# 1  pi=24'b101101110011100000100000;
#1 $display("%b", po);
# 1  pi=24'b101111001101111101111010;
#1 $display("%b", po);
# 1  pi=24'b100110111000110110101001;
#1 $display("%b", po);
# 1  pi=24'b110101001000100101100010;
#1 $display("%b", po);
# 1  pi=24'b011100101000000011011000;
#1 $display("%b", po);
# 1  pi=24'b101001000000000001110000;
#1 $display("%b", po);
# 1  pi=24'b101110110010000100010100;
#1 $display("%b", po);
# 1  pi=24'b011110011000100001100100;
#1 $display("%b", po);
# 1  pi=24'b001100001001110010011010;
#1 $display("%b", po);
# 1  pi=24'b000010010100001010001100;
#1 $display("%b", po);
# 1  pi=24'b101101010101111011101000;
#1 $display("%b", po);
# 1  pi=24'b010111011100110101111001;
#1 $display("%b", po);
# 1  pi=24'b000010100110001110111111;
#1 $display("%b", po);
# 1  pi=24'b000011000100111001110011;
#1 $display("%b", po);
# 1  pi=24'b101100000001100110101011;
#1 $display("%b", po);
# 1  pi=24'b001100011001000010100001;
#1 $display("%b", po);
# 1  pi=24'b101100000011001011000100;
#1 $display("%b", po);
# 1  pi=24'b000001111010101101110010;
#1 $display("%b", po);
# 1  pi=24'b010001001001011000001011;
#1 $display("%b", po);
# 1  pi=24'b010111110111111111011011;
#1 $display("%b", po);
# 1  pi=24'b000000011001001101000000;
#1 $display("%b", po);
# 1  pi=24'b101111000100111111101000;
#1 $display("%b", po);
# 1  pi=24'b110101110111110011100010;
#1 $display("%b", po);
# 1  pi=24'b100000000010100000010000;
#1 $display("%b", po);
# 1  pi=24'b111110111001011000001010;
#1 $display("%b", po);
# 1  pi=24'b100110110101100011101100;
#1 $display("%b", po);
# 1  pi=24'b011101111011011001000000;
#1 $display("%b", po);
# 1  pi=24'b011001011100010001001001;
#1 $display("%b", po);
# 1  pi=24'b011101111101110111101101;
#1 $display("%b", po);
# 1  pi=24'b010111110101001011100110;
#1 $display("%b", po);
# 1  pi=24'b010010011010110111000110;
#1 $display("%b", po);
# 1  pi=24'b111100101000111110110000;
#1 $display("%b", po);
# 1  pi=24'b001100111011100101010100;
#1 $display("%b", po);
# 1  pi=24'b101010010100101000111011;
#1 $display("%b", po);
# 1  pi=24'b001100100111010100100110;
#1 $display("%b", po);
# 1  pi=24'b001111100100110010110010;
#1 $display("%b", po);
# 1  pi=24'b100000100100110010011010;
#1 $display("%b", po);
# 1  pi=24'b001001111101100001101001;
#1 $display("%b", po);
# 1  pi=24'b101011101110000111101010;
#1 $display("%b", po);
# 1  pi=24'b000000101111101101101010;
#1 $display("%b", po);
# 1  pi=24'b010101101110000110100101;
#1 $display("%b", po);
# 1  pi=24'b100111010111000000110010;
#1 $display("%b", po);
# 1  pi=24'b001101011001011001010101;
#1 $display("%b", po);
# 1  pi=24'b000001000110100001011110;
#1 $display("%b", po);
# 1  pi=24'b111000100011010001111011;
#1 $display("%b", po);
# 1  pi=24'b000100110101111110110101;
#1 $display("%b", po);
# 1  pi=24'b001100110000101111110110;
#1 $display("%b", po);
# 1  pi=24'b011111100011011010111001;
#1 $display("%b", po);
# 1  pi=24'b110000111000010010110001;
#1 $display("%b", po);
# 1  pi=24'b011111110000110000001111;
#1 $display("%b", po);
# 1  pi=24'b101111101010110011010001;
#1 $display("%b", po);
# 1  pi=24'b101010110010111001001000;
#1 $display("%b", po);
# 1  pi=24'b100110010111001000111010;
#1 $display("%b", po);
# 1  pi=24'b100110000110011011011101;
#1 $display("%b", po);
# 1  pi=24'b000110110001011000011110;
#1 $display("%b", po);
# 1  pi=24'b011011000001111011000011;
#1 $display("%b", po);
# 1  pi=24'b110010000000100001111011;
#1 $display("%b", po);
# 1  pi=24'b011000001000100110110001;
#1 $display("%b", po);
# 1  pi=24'b100110001101111011001011;
#1 $display("%b", po);
# 1  pi=24'b100000111100110000111010;
#1 $display("%b", po);
# 1  pi=24'b101110101101011100101010;
#1 $display("%b", po);
# 1  pi=24'b011110000011000010000000;
#1 $display("%b", po);
# 1  pi=24'b110010001100000111000111;
#1 $display("%b", po);
# 1  pi=24'b101111111000100011101000;
#1 $display("%b", po);
# 1  pi=24'b001011001100001010100001;
#1 $display("%b", po);
# 1  pi=24'b100100001101100100100100;
#1 $display("%b", po);
# 1  pi=24'b001100111010101101110100;
#1 $display("%b", po);
# 1  pi=24'b010000101101101010101101;
#1 $display("%b", po);
# 1  pi=24'b000011111011010010011100;
#1 $display("%b", po);
# 1  pi=24'b010010111011101110010011;
#1 $display("%b", po);
# 1  pi=24'b100011111101110000100110;
#1 $display("%b", po);
# 1  pi=24'b011011000111011001000010;
#1 $display("%b", po);
# 1  pi=24'b111000101011000000110001;
#1 $display("%b", po);
# 1  pi=24'b010110010001111110011010;
#1 $display("%b", po);
# 1  pi=24'b111010100100110100000101;
#1 $display("%b", po);
# 1  pi=24'b110000111110011000100111;
#1 $display("%b", po);
# 1  pi=24'b111010010110111101000100;
#1 $display("%b", po);
# 1  pi=24'b100100000000010110011100;
#1 $display("%b", po);
# 1  pi=24'b111100101011111110110000;
#1 $display("%b", po);
# 1  pi=24'b010000010010110010101101;
#1 $display("%b", po);
# 1  pi=24'b111110000011001011110111;
#1 $display("%b", po);
# 1  pi=24'b001001001001001010000111;
#1 $display("%b", po);
# 1  pi=24'b001100000100001001100011;
#1 $display("%b", po);
# 1  pi=24'b100100001101111101010111;
#1 $display("%b", po);
# 1  pi=24'b100110000000100101000000;
#1 $display("%b", po);
# 1  pi=24'b001011110000110100000111;
#1 $display("%b", po);
# 1  pi=24'b010111010101011101111110;
#1 $display("%b", po);
# 1  pi=24'b011000110000000000010111;
#1 $display("%b", po);
# 1  pi=24'b111110010001110111011011;
#1 $display("%b", po);
# 1  pi=24'b001001111100111111011110;
#1 $display("%b", po);
# 1  pi=24'b111000010111011101010010;
#1 $display("%b", po);
# 1  pi=24'b111000011001110101101011;
#1 $display("%b", po);
# 1  pi=24'b110111000101000000101110;
#1 $display("%b", po);
# 1  pi=24'b110100111010100010101100;
#1 $display("%b", po);
# 1  pi=24'b010001111010011011110010;
#1 $display("%b", po);
# 1  pi=24'b101001111101101011110010;
#1 $display("%b", po);
# 1  pi=24'b001100111111001011000111;
#1 $display("%b", po);
# 1  pi=24'b110010101000011101010100;
#1 $display("%b", po);
# 1  pi=24'b111111100011101010000111;
#1 $display("%b", po);
# 1  pi=24'b001101000101011101010010;
#1 $display("%b", po);
# 1  pi=24'b101011000001011100001001;
#1 $display("%b", po);
# 1  pi=24'b101011101010111110101011;
#1 $display("%b", po);
# 1  pi=24'b010011010110011100111101;
#1 $display("%b", po);
# 1  pi=24'b000001000000001010001000;
#1 $display("%b", po);
# 1  pi=24'b000001010010001000100010;
#1 $display("%b", po);
# 1  pi=24'b010101011100010011101100;
#1 $display("%b", po);
# 1  pi=24'b100100100011111111010001;
#1 $display("%b", po);
# 1  pi=24'b010001010000000101111111;
#1 $display("%b", po);
# 1  pi=24'b001101000010100100100000;
#1 $display("%b", po);
# 1  pi=24'b001000001001111101101001;
#1 $display("%b", po);
# 1  pi=24'b100010001011011101010000;
#1 $display("%b", po);
# 1  pi=24'b001010101000001111010100;
#1 $display("%b", po);
# 1  pi=24'b010100001000010011001100;
#1 $display("%b", po);
# 1  pi=24'b011111001111000010100011;
#1 $display("%b", po);
# 1  pi=24'b110000011011111010001011;
#1 $display("%b", po);
# 1  pi=24'b101001001010110111010110;
#1 $display("%b", po);
# 1  pi=24'b010100000100110101111000;
#1 $display("%b", po);
# 1  pi=24'b110101000010010110011110;
#1 $display("%b", po);
# 1  pi=24'b011010010010001100001001;
#1 $display("%b", po);
# 1  pi=24'b100110101011111011100011;
#1 $display("%b", po);
# 1  pi=24'b111001101011111100011101;
#1 $display("%b", po);
# 1  pi=24'b010110010001101111111010;
#1 $display("%b", po);
# 1  pi=24'b011100110100101111100100;
#1 $display("%b", po);
# 1  pi=24'b000001010010011101111111;
#1 $display("%b", po);
# 1  pi=24'b010000001011110010111110;
#1 $display("%b", po);
# 1  pi=24'b110110001000010101000111;
#1 $display("%b", po);
# 1  pi=24'b111011011111100011110110;
#1 $display("%b", po);
# 1  pi=24'b010111000101001101001110;
#1 $display("%b", po);
# 1  pi=24'b111110010110011010001010;
#1 $display("%b", po);
# 1  pi=24'b110000000111010110100110;
#1 $display("%b", po);
# 1  pi=24'b100001011001101100110000;
#1 $display("%b", po);
# 1  pi=24'b110001011110100000100011;
#1 $display("%b", po);
# 1  pi=24'b010011001010010101110100;
#1 $display("%b", po);
# 1  pi=24'b011001101011111010111110;
#1 $display("%b", po);
# 1  pi=24'b101011111010101101100110;
#1 $display("%b", po);
# 1  pi=24'b101110000110010110000100;
#1 $display("%b", po);
# 1  pi=24'b000101111100111111000101;
#1 $display("%b", po);
# 1  pi=24'b011000000010101111100000;
#1 $display("%b", po);
# 1  pi=24'b001011010011010011010111;
#1 $display("%b", po);
# 1  pi=24'b101000100101000100010001;
#1 $display("%b", po);
# 1  pi=24'b111110010011010000011011;
#1 $display("%b", po);
# 1  pi=24'b111100011001010000000011;
#1 $display("%b", po);
# 1  pi=24'b101100010000110110111111;
#1 $display("%b", po);
# 1  pi=24'b000111101001000011000000;
#1 $display("%b", po);
# 1  pi=24'b000111110101010001101101;
#1 $display("%b", po);
# 1  pi=24'b001111101100111100010001;
#1 $display("%b", po);
# 1  pi=24'b110110010100001000000000;
#1 $display("%b", po);
# 1  pi=24'b111011101001101101000101;
#1 $display("%b", po);
# 1  pi=24'b101010110110100111010110;
#1 $display("%b", po);
# 1  pi=24'b000100010010000010101101;
#1 $display("%b", po);
# 1  pi=24'b000110110110110010110111;
#1 $display("%b", po);
# 1  pi=24'b110000011010000000011110;
#1 $display("%b", po);
# 1  pi=24'b000011001111111100001010;
#1 $display("%b", po);
# 1  pi=24'b001010001110101001010101;
#1 $display("%b", po);
# 1  pi=24'b010001000101110100011111;
#1 $display("%b", po);
# 1  pi=24'b111110000010011111001101;
#1 $display("%b", po);
# 1  pi=24'b011101010010010101100100;
#1 $display("%b", po);
# 1  pi=24'b100101011111111110110100;
#1 $display("%b", po);
# 1  pi=24'b100111110001011100001100;
#1 $display("%b", po);
# 1  pi=24'b000010101010000011001100;
#1 $display("%b", po);
# 1  pi=24'b011011110001110101101001;
#1 $display("%b", po);
# 1  pi=24'b011101101101000110011001;
#1 $display("%b", po);
# 1  pi=24'b110011101111110100001010;
#1 $display("%b", po);
# 1  pi=24'b100000101110110110101111;
#1 $display("%b", po);
# 1  pi=24'b011001010001000101100100;
#1 $display("%b", po);
# 1  pi=24'b000110000011101010011001;
#1 $display("%b", po);
# 1  pi=24'b101001001110110010100010;
#1 $display("%b", po);
# 1  pi=24'b010010000100100101110000;
#1 $display("%b", po);
# 1  pi=24'b011011001011100101001010;
#1 $display("%b", po);
# 1  pi=24'b011111010110011111110100;
#1 $display("%b", po);
# 1  pi=24'b000001011100100100010000;
#1 $display("%b", po);
# 1  pi=24'b010001011001001001001001;
#1 $display("%b", po);
# 1  pi=24'b011100011000100011000010;
#1 $display("%b", po);
# 1  pi=24'b100111000010011100110110;
#1 $display("%b", po);
# 1  pi=24'b000000111100001000001110;
#1 $display("%b", po);
# 1  pi=24'b101000101010011010000101;
#1 $display("%b", po);
# 1  pi=24'b001001011000000011010111;
#1 $display("%b", po);
# 1  pi=24'b111111110111001111101101;
#1 $display("%b", po);
# 1  pi=24'b100100111111010001001011;
#1 $display("%b", po);
# 1  pi=24'b100010111001000011111001;
#1 $display("%b", po);
# 1  pi=24'b101010011011101111011011;
#1 $display("%b", po);
# 1  pi=24'b101011000100001000010011;
#1 $display("%b", po);
# 1  pi=24'b011000001111100001111100;
#1 $display("%b", po);
# 1  pi=24'b011110001110110100000100;
#1 $display("%b", po);
# 1  pi=24'b000000011101000010100101;
#1 $display("%b", po);
# 1  pi=24'b010001101011011000001101;
#1 $display("%b", po);
# 1  pi=24'b000011100011110011100101;
#1 $display("%b", po);
# 1  pi=24'b010000100110110000001111;
#1 $display("%b", po);
# 1  pi=24'b001011011011010111011111;
#1 $display("%b", po);
# 1  pi=24'b001000111000001010111100;
#1 $display("%b", po);
# 1  pi=24'b010110110110011001000000;
#1 $display("%b", po);
# 1  pi=24'b011101100001110011011100;
#1 $display("%b", po);
# 1  pi=24'b110101010111110111110011;
#1 $display("%b", po);
# 1  pi=24'b111001101001011000011101;
#1 $display("%b", po);
# 1  pi=24'b110011110011000011111011;
#1 $display("%b", po);
# 1  pi=24'b110100110010001011101000;
#1 $display("%b", po);
# 1  pi=24'b100110110100101000000011;
#1 $display("%b", po);
# 1  pi=24'b001101111001010011010011;
#1 $display("%b", po);
# 1  pi=24'b110011010010011100111010;
#1 $display("%b", po);
# 1  pi=24'b001100100011011100100010;
#1 $display("%b", po);
# 1  pi=24'b111111001001011111010001;
#1 $display("%b", po);
# 1  pi=24'b100011101110101110111101;
#1 $display("%b", po);
# 1  pi=24'b000111111000100010101101;
#1 $display("%b", po);
# 1  pi=24'b100010010100001011111100;
#1 $display("%b", po);
# 1  pi=24'b110100100111001001110100;
#1 $display("%b", po);
# 1  pi=24'b011000010101100011000010;
#1 $display("%b", po);
# 1  pi=24'b101001100001010111011100;
#1 $display("%b", po);
# 1  pi=24'b000110100001110110001010;
#1 $display("%b", po);
# 1  pi=24'b111001111001101101111101;
#1 $display("%b", po);
# 1  pi=24'b001101110010011110011011;
#1 $display("%b", po);
# 1  pi=24'b101011110111111110010011;
#1 $display("%b", po);
# 1  pi=24'b000101111100010101100010;
#1 $display("%b", po);
# 1  pi=24'b011101101000101100101000;
#1 $display("%b", po);
# 1  pi=24'b100000110001000000001000;
#1 $display("%b", po);
# 1  pi=24'b110100111101010100001010;
#1 $display("%b", po);
# 1  pi=24'b110100000100110111011111;
#1 $display("%b", po);
# 1  pi=24'b010010110000010001000101;
#1 $display("%b", po);
# 1  pi=24'b010110111001100110100011;
#1 $display("%b", po);
# 1  pi=24'b101010000010000110000010;
#1 $display("%b", po);
# 1  pi=24'b111001101010000110011001;
#1 $display("%b", po);
# 1  pi=24'b101101001101100000100001;
#1 $display("%b", po);
# 1  pi=24'b001101001010010111100111;
#1 $display("%b", po);
# 1  pi=24'b011110011101000011001000;
#1 $display("%b", po);
# 1  pi=24'b000111010010101100001001;
#1 $display("%b", po);
# 1  pi=24'b110111111100100111001100;
#1 $display("%b", po);
# 1  pi=24'b100111000000101000001111;
#1 $display("%b", po);
# 1  pi=24'b100011011111110101010000;
#1 $display("%b", po);
# 1  pi=24'b010010001001111110001010;
#1 $display("%b", po);
# 1  pi=24'b000001110011010111111111;
#1 $display("%b", po);
# 1  pi=24'b111001000000110101000110;
#1 $display("%b", po);
# 1  pi=24'b001010011110001000001000;
#1 $display("%b", po);
# 1  pi=24'b110111000111110101101111;
#1 $display("%b", po);
# 1  pi=24'b110111010100001110100100;
#1 $display("%b", po);
# 1  pi=24'b100011101001001100010110;
#1 $display("%b", po);
# 1  pi=24'b100100111111110001010100;
#1 $display("%b", po);
# 1  pi=24'b111100000000101111000101;
#1 $display("%b", po);
# 1  pi=24'b111000000101111001110101;
#1 $display("%b", po);
# 1  pi=24'b101000111010001101101000;
#1 $display("%b", po);
# 1  pi=24'b010001011111111110011010;
#1 $display("%b", po);
# 1  pi=24'b100000110111111001101010;
#1 $display("%b", po);
# 1  pi=24'b011101001101101110010011;
#1 $display("%b", po);
# 1  pi=24'b010010100101101110100101;
#1 $display("%b", po);
# 1  pi=24'b111101101110111101110001;
#1 $display("%b", po);
# 1  pi=24'b011001000010010010001110;
#1 $display("%b", po);
# 1  pi=24'b000001010110011100111111;
#1 $display("%b", po);
# 1  pi=24'b010010101011110000000110;
#1 $display("%b", po);
# 1  pi=24'b011000101010110101100011;
#1 $display("%b", po);
# 1  pi=24'b010100011011001111110100;
#1 $display("%b", po);
# 1  pi=24'b100000111110001101101000;
#1 $display("%b", po);
# 1  pi=24'b010111000110001010011000;
#1 $display("%b", po);
# 1  pi=24'b010100011100101010011010;
#1 $display("%b", po);
# 1  pi=24'b111000110001100110011000;
#1 $display("%b", po);
# 1  pi=24'b010011111110100101011001;
#1 $display("%b", po);
# 1  pi=24'b111010011110000000001000;
#1 $display("%b", po);
# 1  pi=24'b000110000111100010100001;
#1 $display("%b", po);
# 1  pi=24'b101110011001110010001010;
#1 $display("%b", po);
# 1  pi=24'b001011111110010010011001;
#1 $display("%b", po);
# 1  pi=24'b100001001010010011110000;
#1 $display("%b", po);
# 1  pi=24'b100101011000100010101000;
#1 $display("%b", po);
# 1  pi=24'b011011110101111010000000;
#1 $display("%b", po);
# 1  pi=24'b001000010110110101100011;
#1 $display("%b", po);
# 1  pi=24'b000000111111010111110011;
#1 $display("%b", po);
# 1  pi=24'b001000010000110100110011;
#1 $display("%b", po);
# 1  pi=24'b010101010000101011110001;
#1 $display("%b", po);
# 1  pi=24'b010000010011010011010100;
#1 $display("%b", po);
# 1  pi=24'b000011100001110011011100;
#1 $display("%b", po);
# 1  pi=24'b100101000100101010110100;
#1 $display("%b", po);
# 1  pi=24'b001111010000000110100111;
#1 $display("%b", po);
# 1  pi=24'b101101011010100111011100;
#1 $display("%b", po);
# 1  pi=24'b001010100101110100101001;
#1 $display("%b", po);
# 1  pi=24'b110110100111110101000010;
#1 $display("%b", po);
# 1  pi=24'b000111100111010101000001;
#1 $display("%b", po);
# 1  pi=24'b011111001101010001110011;
#1 $display("%b", po);
# 1  pi=24'b100100100010110000011111;
#1 $display("%b", po);
# 1  pi=24'b000100011101011110011110;
#1 $display("%b", po);
# 1  pi=24'b011000010101010111111111;
#1 $display("%b", po);
# 1  pi=24'b110110111001110001010110;
#1 $display("%b", po);
# 1  pi=24'b101100110011101000000001;
#1 $display("%b", po);
# 1  pi=24'b110001101000000100101111;
#1 $display("%b", po);
# 1  pi=24'b001101001101011000000100;
#1 $display("%b", po);
# 1  pi=24'b100110110110000010100011;
#1 $display("%b", po);
# 1  pi=24'b011010000101011001001010;
#1 $display("%b", po);
# 1  pi=24'b000011101001101011001010;
#1 $display("%b", po);
# 1  pi=24'b000000111101000011101001;
#1 $display("%b", po);
# 1  pi=24'b011110011011100110100000;
#1 $display("%b", po);
# 1  pi=24'b001010111111001010001110;
#1 $display("%b", po);
# 1  pi=24'b111010001001001011110101;
#1 $display("%b", po);
# 1  pi=24'b101001010110101100001010;
#1 $display("%b", po);
# 1  pi=24'b101011011101100101100000;
#1 $display("%b", po);
# 1  pi=24'b000110101011111101011010;
#1 $display("%b", po);
# 1  pi=24'b110100110111100000011101;
#1 $display("%b", po);
# 1  pi=24'b101110111011101001011011;
#1 $display("%b", po);
# 1  pi=24'b010001001011011010010100;
#1 $display("%b", po);
# 1  pi=24'b111111100010001100101000;
#1 $display("%b", po);
# 1  pi=24'b011101101101010011011100;
#1 $display("%b", po);
# 1  pi=24'b100011011001001010111110;
#1 $display("%b", po);
# 1  pi=24'b100000001111101110011001;
#1 $display("%b", po);
# 1  pi=24'b010111111011101011101000;
#1 $display("%b", po);
# 1  pi=24'b001110010101001100010000;
#1 $display("%b", po);
# 1  pi=24'b110100010001110010111111;
#1 $display("%b", po);
# 1  pi=24'b010101001001110100101000;
#1 $display("%b", po);
# 1  pi=24'b111101010101111000111101;
#1 $display("%b", po);
# 1  pi=24'b010100111010011000000000;
#1 $display("%b", po);
# 1  pi=24'b111000111101001110100100;
#1 $display("%b", po);
# 1  pi=24'b011101110100111001010111;
#1 $display("%b", po);
# 1  pi=24'b111101000110100101011111;
#1 $display("%b", po);
# 1  pi=24'b000100100101101001101011;
#1 $display("%b", po);
# 1  pi=24'b000101110110100111010011;
#1 $display("%b", po);
# 1  pi=24'b000000011111111010100101;
#1 $display("%b", po);
# 1  pi=24'b001010110100000100000101;
#1 $display("%b", po);
# 1  pi=24'b101000111101110001101011;
#1 $display("%b", po);
# 1  pi=24'b100010100111110100110111;
#1 $display("%b", po);
# 1  pi=24'b100100110011110101100011;
#1 $display("%b", po);
# 1  pi=24'b011000001110010001010100;
#1 $display("%b", po);
# 1  pi=24'b001110000010110101111111;
#1 $display("%b", po);
# 1  pi=24'b111000010111001000010111;
#1 $display("%b", po);
# 1  pi=24'b000100010010011000001001;
#1 $display("%b", po);
# 1  pi=24'b110110111000100110011011;
#1 $display("%b", po);
# 1  pi=24'b011101000111011101001011;
#1 $display("%b", po);
# 1  pi=24'b000100001110101100101001;
#1 $display("%b", po);
# 1  pi=24'b101011000010100111100011;
#1 $display("%b", po);
# 1  pi=24'b100110010110111011110111;
#1 $display("%b", po);
# 1  pi=24'b001110100001001011010110;
#1 $display("%b", po);
# 1  pi=24'b101101011110011001010101;
#1 $display("%b", po);
# 1  pi=24'b011011100111011101010110;
#1 $display("%b", po);
# 1  pi=24'b000000110000010011000111;
#1 $display("%b", po);
# 1  pi=24'b110011101101101000011110;
#1 $display("%b", po);
# 1  pi=24'b010001001010101010110110;
#1 $display("%b", po);
# 1  pi=24'b111100010011111110101101;
#1 $display("%b", po);
# 1  pi=24'b010111011101101111111101;
#1 $display("%b", po);
# 1  pi=24'b010000111111101110110001;
#1 $display("%b", po);
# 1  pi=24'b010100000111011010100110;
#1 $display("%b", po);
# 1  pi=24'b010001111111101010001110;
#1 $display("%b", po);
# 1  pi=24'b000000111110001000110101;
#1 $display("%b", po);
# 1  pi=24'b111000110001000001100010;
#1 $display("%b", po);
# 1  pi=24'b111110111000010011000011;
#1 $display("%b", po);
# 1  pi=24'b011000001100000010110001;
#1 $display("%b", po);
# 1  pi=24'b101110010001100101001011;
#1 $display("%b", po);
# 1  pi=24'b000100000110110100100100;
#1 $display("%b", po);
# 1  pi=24'b001110011111100100000110;
#1 $display("%b", po);
# 1  pi=24'b011101100101110000001100;
#1 $display("%b", po);
# 1  pi=24'b001101001011110110111100;
#1 $display("%b", po);
# 1  pi=24'b100101100111000001011100;
#1 $display("%b", po);
# 1  pi=24'b001111111001110100100111;
#1 $display("%b", po);
# 1  pi=24'b001010100111101100000100;
#1 $display("%b", po);
# 1  pi=24'b101010011101110010111011;
#1 $display("%b", po);
# 1  pi=24'b100101000110101011101110;
#1 $display("%b", po);
# 1  pi=24'b111110110001111100101010;
#1 $display("%b", po);
# 1  pi=24'b011011101011110111011111;
#1 $display("%b", po);
# 1  pi=24'b110101010110011111001010;
#1 $display("%b", po);
# 1  pi=24'b110111001111011001101010;
#1 $display("%b", po);
# 1  pi=24'b111000100110111110101001;
#1 $display("%b", po);
# 1  pi=24'b111100010110111011010001;
#1 $display("%b", po);
# 1  pi=24'b101011010100000001110110;
#1 $display("%b", po);
# 1  pi=24'b111100001111011010100010;
#1 $display("%b", po);
# 1  pi=24'b101000011110001110110110;
#1 $display("%b", po);
# 1  pi=24'b100110111010110110010101;
#1 $display("%b", po);
# 1  pi=24'b000001111001000011001111;
#1 $display("%b", po);
# 1  pi=24'b110000001000110110010010;
#1 $display("%b", po);
# 1  pi=24'b111010100101011000010111;
#1 $display("%b", po);
# 1  pi=24'b001101100000010000010110;
#1 $display("%b", po);
# 1  pi=24'b011110001110000011010011;
#1 $display("%b", po);
# 1  pi=24'b000111010111111100100000;
#1 $display("%b", po);
# 1  pi=24'b111001001100001110011101;
#1 $display("%b", po);
# 1  pi=24'b101101101101101100001001;
#1 $display("%b", po);
# 1  pi=24'b010100010101100110010011;
#1 $display("%b", po);
# 1  pi=24'b011000001100111111011111;
#1 $display("%b", po);
# 1  pi=24'b111011100001100001000011;
#1 $display("%b", po);
# 1  pi=24'b011100010100100010110011;
#1 $display("%b", po);
# 1  pi=24'b011100100011000011011110;
#1 $display("%b", po);
# 1  pi=24'b001101000001001100110001;
#1 $display("%b", po);
# 1  pi=24'b000111111001101011111011;
#1 $display("%b", po);
# 1  pi=24'b001110010100111101010001;
#1 $display("%b", po);
# 1  pi=24'b001001001100000110101000;
#1 $display("%b", po);
# 1  pi=24'b010000100110000010110011;
#1 $display("%b", po);
# 1  pi=24'b000001101011100001100101;
#1 $display("%b", po);
# 1  pi=24'b100000011001110000010110;
#1 $display("%b", po);
# 1  pi=24'b001111101111010111101001;
#1 $display("%b", po);
# 1  pi=24'b100100000010111010101111;
#1 $display("%b", po);
# 1  pi=24'b111110110001111100110000;
#1 $display("%b", po);
# 1  pi=24'b000000000100011111111101;
#1 $display("%b", po);
# 1  pi=24'b110001110100000010110110;
#1 $display("%b", po);
# 1  pi=24'b011111101001000110000010;
#1 $display("%b", po);
# 1  pi=24'b000111000011110100001111;
#1 $display("%b", po);
# 1  pi=24'b111000010011100100101010;
#1 $display("%b", po);
# 1  pi=24'b101100000110000010100110;
#1 $display("%b", po);
# 1  pi=24'b110110110100001110011011;
#1 $display("%b", po);
# 1  pi=24'b100001001111111101111101;
#1 $display("%b", po);
# 1  pi=24'b110111011101110101101001;
#1 $display("%b", po);
# 1  pi=24'b001100000001010010011000;
#1 $display("%b", po);
# 1  pi=24'b110101011111100111011001;
#1 $display("%b", po);
# 1  pi=24'b001001010011101111001010;
#1 $display("%b", po);
# 1  pi=24'b110101111001001011010000;
#1 $display("%b", po);
# 1  pi=24'b100001011100100000000011;
#1 $display("%b", po);
# 1  pi=24'b001010001010001100100001;
#1 $display("%b", po);
# 1  pi=24'b010100100000101001110111;
#1 $display("%b", po);
# 1  pi=24'b100111111001111110111000;
#1 $display("%b", po);
# 1  pi=24'b001111111010110001110011;
#1 $display("%b", po);
# 1  pi=24'b100010001011011100110010;
#1 $display("%b", po);
# 1  pi=24'b101100101101100000110111;
#1 $display("%b", po);
# 1  pi=24'b010110111011011011000101;
#1 $display("%b", po);
# 1  pi=24'b001110000100010001100000;
#1 $display("%b", po);
# 1  pi=24'b010111100001100001001111;
#1 $display("%b", po);
# 1  pi=24'b010010000010000000111010;
#1 $display("%b", po);
# 1  pi=24'b100111010111101111000010;
#1 $display("%b", po);
# 1  pi=24'b000100110001101001110100;
#1 $display("%b", po);
# 1  pi=24'b101001111010100010101010;
#1 $display("%b", po);
# 1  pi=24'b000010110001111111000101;
#1 $display("%b", po);
# 1  pi=24'b000101011110001100111110;
#1 $display("%b", po);
# 1  pi=24'b010010010110101011001001;
#1 $display("%b", po);
# 1  pi=24'b100111001111111010110011;
#1 $display("%b", po);
# 1  pi=24'b001110101001000001111001;
#1 $display("%b", po);
# 1  pi=24'b010110011100011001000010;
#1 $display("%b", po);
# 1  pi=24'b000111111001001010001111;
#1 $display("%b", po);
# 1  pi=24'b010000101101000111001000;
#1 $display("%b", po);
# 1  pi=24'b100111110000110011010101;
#1 $display("%b", po);
# 1  pi=24'b101110001000110010111100;
#1 $display("%b", po);
# 1  pi=24'b111001111010000010111101;
#1 $display("%b", po);
# 1  pi=24'b110110000110101100001101;
#1 $display("%b", po);
# 1  pi=24'b110001101111100111010111;
#1 $display("%b", po);
# 1  pi=24'b101110100010011110001001;
#1 $display("%b", po);
# 1  pi=24'b000110101100110000110010;
#1 $display("%b", po);
# 1  pi=24'b101101010101001010000011;
#1 $display("%b", po);
# 1  pi=24'b111111100111000011010111;
#1 $display("%b", po);
# 1  pi=24'b110001000111001100110011;
#1 $display("%b", po);
# 1  pi=24'b011011001101101111011010;
#1 $display("%b", po);
# 1  pi=24'b101111000000100110111001;
#1 $display("%b", po);
# 1  pi=24'b010011110010100011010111;
#1 $display("%b", po);
# 1  pi=24'b000111111101110101111000;
#1 $display("%b", po);
# 1  pi=24'b111111111100000011100011;
#1 $display("%b", po);
# 1  pi=24'b001101110000010011101110;
#1 $display("%b", po);
# 1  pi=24'b011010010001000110001110;
#1 $display("%b", po);
# 1  pi=24'b101100011101000111100001;
#1 $display("%b", po);
# 1  pi=24'b100101101100101101101011;
#1 $display("%b", po);
# 1  pi=24'b101111110001110001010000;
#1 $display("%b", po);
# 1  pi=24'b011101111101111000011111;
#1 $display("%b", po);
# 1  pi=24'b001101110101011001111000;
#1 $display("%b", po);
# 1  pi=24'b110010000111111111000011;
#1 $display("%b", po);
# 1  pi=24'b100011010010100111010101;
#1 $display("%b", po);
# 1  pi=24'b010001001111010001010110;
#1 $display("%b", po);
# 1  pi=24'b011001100111011100010000;
#1 $display("%b", po);
# 1  pi=24'b111010111000010100001111;
#1 $display("%b", po);
# 1  pi=24'b011110110110110101110011;
#1 $display("%b", po);
# 1  pi=24'b001100011010111100100100;
#1 $display("%b", po);
# 1  pi=24'b110011111011001110001100;
#1 $display("%b", po);
# 1  pi=24'b100101001111010000110101;
#1 $display("%b", po);
# 1  pi=24'b001001110001100011110110;
#1 $display("%b", po);
# 1  pi=24'b010110001110101000111111;
#1 $display("%b", po);
# 1  pi=24'b101111100001000100110001;
#1 $display("%b", po);
# 1  pi=24'b100110000001111000010101;
#1 $display("%b", po);
# 1  pi=24'b111000001101111100011001;
#1 $display("%b", po);
# 1  pi=24'b000101010010111000110111;
#1 $display("%b", po);
# 1  pi=24'b011101010101010000101100;
#1 $display("%b", po);
# 1  pi=24'b111110001011000111100100;
#1 $display("%b", po);
# 1  pi=24'b001010000001000100000101;
#1 $display("%b", po);
# 1  pi=24'b111111100101011000000111;
#1 $display("%b", po);
# 1  pi=24'b110110101110111010010110;
#1 $display("%b", po);
# 1  pi=24'b000000011111110110011110;
#1 $display("%b", po);
# 1  pi=24'b000100110110000011000100;
#1 $display("%b", po);
# 1  pi=24'b001001010010101000010001;
#1 $display("%b", po);
# 1  pi=24'b101000011001011011101011;
#1 $display("%b", po);
# 1  pi=24'b000011110111111100110111;
#1 $display("%b", po);
# 1  pi=24'b111100101110010000100010;
#1 $display("%b", po);
# 1  pi=24'b110010000010100001100010;
#1 $display("%b", po);
# 1  pi=24'b010101101101100011011010;
#1 $display("%b", po);
# 1  pi=24'b001111111001011101010010;
#1 $display("%b", po);
# 1  pi=24'b011000111010000011111000;
#1 $display("%b", po);
# 1  pi=24'b001001010001010011001111;
#1 $display("%b", po);
# 1  pi=24'b100110101001100000010101;
#1 $display("%b", po);
# 1  pi=24'b100010100000001111101001;
#1 $display("%b", po);
# 1  pi=24'b110001100001001011010111;
#1 $display("%b", po);
# 1  pi=24'b010100000000001111011001;
#1 $display("%b", po);
# 1  pi=24'b110110001111111001100000;
#1 $display("%b", po);
# 1  pi=24'b011101000101000011000100;
#1 $display("%b", po);
# 1  pi=24'b011000001000000010011100;
#1 $display("%b", po);
# 1  pi=24'b010001010000110011000011;
#1 $display("%b", po);
# 1  pi=24'b101011110100111010010000;
#1 $display("%b", po);
# 1  pi=24'b011111000101100001011010;
#1 $display("%b", po);
# 1  pi=24'b001110000000101110100110;
#1 $display("%b", po);
# 1  pi=24'b110110001110000000110101;
#1 $display("%b", po);
# 1  pi=24'b000001001010100101110100;
#1 $display("%b", po);
# 1  pi=24'b000111101011101000101000;
#1 $display("%b", po);
# 1  pi=24'b010110110010010000110001;
#1 $display("%b", po);
# 1  pi=24'b001010000010000010101110;
#1 $display("%b", po);
# 1  pi=24'b010000000110100100000011;
#1 $display("%b", po);
# 1  pi=24'b000010110011101111100010;
#1 $display("%b", po);
# 1  pi=24'b010100010101100101100101;
#1 $display("%b", po);
# 1  pi=24'b011001011010110101011111;
#1 $display("%b", po);
# 1  pi=24'b001001010000101101001011;
#1 $display("%b", po);
# 1  pi=24'b100110100011111110000111;
#1 $display("%b", po);
# 1  pi=24'b010011011010101010000110;
#1 $display("%b", po);
# 1  pi=24'b010101010110011000100111;
#1 $display("%b", po);
# 1  pi=24'b100110010001000100010100;
#1 $display("%b", po);
# 1  pi=24'b101011100110000100011010;
#1 $display("%b", po);
# 1  pi=24'b111001101110010100001101;
#1 $display("%b", po);
# 1  pi=24'b000101111011110101110000;
#1 $display("%b", po);
# 1  pi=24'b010110001011010110101010;
#1 $display("%b", po);
# 1  pi=24'b101111101101000000110100;
#1 $display("%b", po);
# 1  pi=24'b111001010110100100100110;
#1 $display("%b", po);
# 1  pi=24'b010100001110111111010001;
#1 $display("%b", po);
# 1  pi=24'b110011000011000011101010;
#1 $display("%b", po);
# 1  pi=24'b010100100001001101110011;
#1 $display("%b", po);
# 1  pi=24'b110101001011100000011100;
#1 $display("%b", po);
# 1  pi=24'b001111110111111011000001;
#1 $display("%b", po);
# 1  pi=24'b010101010110001111100111;
#1 $display("%b", po);
# 1  pi=24'b110001111110010100001000;
#1 $display("%b", po);
# 1  pi=24'b011101011100001010100111;
#1 $display("%b", po);
# 1  pi=24'b101101010101101110001110;
#1 $display("%b", po);
# 1  pi=24'b000001001111101110000001;
#1 $display("%b", po);
# 1  pi=24'b000010000110111111110001;
#1 $display("%b", po);
# 1  pi=24'b110001100110010010000001;
#1 $display("%b", po);
# 1  pi=24'b000000001110110101100111;
#1 $display("%b", po);
# 1  pi=24'b110101011000001111001011;
#1 $display("%b", po);
# 1  pi=24'b011100000111010011111001;
#1 $display("%b", po);
# 1  pi=24'b000100100011011000111110;
#1 $display("%b", po);
# 1  pi=24'b010011101010000011101011;
#1 $display("%b", po);
# 1  pi=24'b110001011110010001001000;
#1 $display("%b", po);
# 1  pi=24'b101101011000000000101100;
#1 $display("%b", po);
# 1  pi=24'b000111101001111011010111;
#1 $display("%b", po);
# 1  pi=24'b001011000111011111101001;
#1 $display("%b", po);
# 1  pi=24'b110001011100010111011001;
#1 $display("%b", po);
# 1  pi=24'b111011111001111110111001;
#1 $display("%b", po);
# 1  pi=24'b111110011000110100010100;
#1 $display("%b", po);
# 1  pi=24'b001101101010110011010111;
#1 $display("%b", po);
# 1  pi=24'b000100001100010000101010;
#1 $display("%b", po);
# 1  pi=24'b010010100110001011001011;
#1 $display("%b", po);
# 1  pi=24'b101011000011010010101100;
#1 $display("%b", po);
# 1  pi=24'b111110001101111011100001;
#1 $display("%b", po);
# 1  pi=24'b011010000001000111111101;
#1 $display("%b", po);
# 1  pi=24'b011110110111111101101101;
#1 $display("%b", po);
# 1  pi=24'b000101100001111001011111;
#1 $display("%b", po);
# 1  pi=24'b100000001101010110001000;
#1 $display("%b", po);
# 1  pi=24'b101011111000111101000000;
#1 $display("%b", po);
# 1  pi=24'b100111111100001110000101;
#1 $display("%b", po);
# 1  pi=24'b010000101101001100101001;
#1 $display("%b", po);
# 1  pi=24'b011100000001001010101000;
#1 $display("%b", po);
# 1  pi=24'b010110110111100111101100;
#1 $display("%b", po);
# 1  pi=24'b101110001011100001100000;
#1 $display("%b", po);
# 1  pi=24'b100011010100011100001001;
#1 $display("%b", po);
# 1  pi=24'b100110100000110001001000;
#1 $display("%b", po);
# 1  pi=24'b111101000100101110000011;
#1 $display("%b", po);
# 1  pi=24'b010100001000110100100111;
#1 $display("%b", po);
# 1  pi=24'b100000110011111011100000;
#1 $display("%b", po);
# 1  pi=24'b011011100011010001100000;
#1 $display("%b", po);
# 1  pi=24'b111001011100100001111111;
#1 $display("%b", po);
# 1  pi=24'b110111101001010011010011;
#1 $display("%b", po);
# 1  pi=24'b110010000110000101110111;
#1 $display("%b", po);
# 1  pi=24'b111010010100110101001111;
#1 $display("%b", po);
# 1  pi=24'b110100110010000001000001;
#1 $display("%b", po);
# 1  pi=24'b001111000111001010011110;
#1 $display("%b", po);
# 1  pi=24'b011100000001000010011100;
#1 $display("%b", po);
# 1  pi=24'b000000010011011000110101;
#1 $display("%b", po);
# 1  pi=24'b101101111011000100111110;
#1 $display("%b", po);
# 1  pi=24'b001000001001110111100110;
#1 $display("%b", po);
# 1  pi=24'b010010001100000100010010;
#1 $display("%b", po);
# 1  pi=24'b000010101010000001001101;
#1 $display("%b", po);
# 1  pi=24'b000010100111100100100001;
#1 $display("%b", po);
# 1  pi=24'b011001001100001101101001;
#1 $display("%b", po);
# 1  pi=24'b110101010011000000001011;
#1 $display("%b", po);
# 1  pi=24'b011000011011010110100010;
#1 $display("%b", po);
# 1  pi=24'b111011101000010100110001;
#1 $display("%b", po);
# 1  pi=24'b001000101001000010001100;
#1 $display("%b", po);
# 1  pi=24'b001011100010010101101001;
#1 $display("%b", po);
# 1  pi=24'b001110110011011000000100;
#1 $display("%b", po);
# 1  pi=24'b111001001110001100010111;
#1 $display("%b", po);
# 1  pi=24'b100111110011101001001100;
#1 $display("%b", po);
# 1  pi=24'b101010101001101011000001;
#1 $display("%b", po);
# 1  pi=24'b100001110100000011011110;
#1 $display("%b", po);
# 1  pi=24'b111101010001100011001111;
#1 $display("%b", po);
# 1  pi=24'b111111101110100000101111;
#1 $display("%b", po);
# 1  pi=24'b101010110010110001111000;
#1 $display("%b", po);
# 1  pi=24'b001100111100001100111100;
#1 $display("%b", po);
# 1  pi=24'b000111001000101111000010;
#1 $display("%b", po);
# 1  pi=24'b101000010000111100010111;
#1 $display("%b", po);
# 1  pi=24'b100001010000101110101100;
#1 $display("%b", po);
# 1  pi=24'b001111010001001101010011;
#1 $display("%b", po);
# 1  pi=24'b011101100101000100010111;
#1 $display("%b", po);
# 1  pi=24'b110111011011111010011100;
#1 $display("%b", po);
# 1  pi=24'b110000110100010110001010;
#1 $display("%b", po);
# 1  pi=24'b001111111000111011111001;
#1 $display("%b", po);
# 1  pi=24'b111001000000000001010001;
#1 $display("%b", po);
# 1  pi=24'b100011000000101111010001;
#1 $display("%b", po);
# 1  pi=24'b100010100111100110001010;
#1 $display("%b", po);
# 1  pi=24'b110010011101001011111011;
#1 $display("%b", po);
# 1  pi=24'b100110111011100111110101;
#1 $display("%b", po);
# 1  pi=24'b111101101000101111101010;
#1 $display("%b", po);
# 1  pi=24'b110011101101110100101011;
#1 $display("%b", po);
# 1  pi=24'b011101111100000111001101;
#1 $display("%b", po);
# 1  pi=24'b010110110010100000101011;
#1 $display("%b", po);
# 1  pi=24'b001011110011101110101001;
#1 $display("%b", po);
# 1  pi=24'b000101010000100110011100;
#1 $display("%b", po);
# 1  pi=24'b110011111011101011000110;
#1 $display("%b", po);
# 1  pi=24'b010110011110000110100100;
#1 $display("%b", po);
# 1  pi=24'b011111011100101011000000;
#1 $display("%b", po);
# 1  pi=24'b000001101000010100100000;
#1 $display("%b", po);
# 1  pi=24'b000101101010111001110110;
#1 $display("%b", po);
# 1  pi=24'b010001110011011011000111;
#1 $display("%b", po);
# 1  pi=24'b000010011011001010101011;
#1 $display("%b", po);
# 1  pi=24'b001110100111010000001100;
#1 $display("%b", po);
# 1  pi=24'b011101101000100010111011;
#1 $display("%b", po);
# 1  pi=24'b011111100110111100011101;
#1 $display("%b", po);
# 1  pi=24'b101101101001000111101100;
#1 $display("%b", po);
# 1  pi=24'b101010110100001110011101;
#1 $display("%b", po);
# 1  pi=24'b101011001101101001101010;
#1 $display("%b", po);
# 1  pi=24'b100101011000110111111110;
#1 $display("%b", po);
# 1  pi=24'b111100010111000000101111;
#1 $display("%b", po);
# 1  pi=24'b011011000010010101100000;
#1 $display("%b", po);
# 1  pi=24'b100111011111100000110101;
#1 $display("%b", po);
# 1  pi=24'b101010011101000101100110;
#1 $display("%b", po);
# 1  pi=24'b001100010010011111111100;
#1 $display("%b", po);
# 1  pi=24'b111111101111000001000110;
#1 $display("%b", po);
# 1  pi=24'b000101000101010110010010;
#1 $display("%b", po);
# 1  pi=24'b100111000101010011101010;
#1 $display("%b", po);
# 1  pi=24'b011001000110101011100000;
#1 $display("%b", po);
# 1  pi=24'b011011101101011101100011;
#1 $display("%b", po);
# 1  pi=24'b001011101110000011000110;
#1 $display("%b", po);
# 1  pi=24'b110010101100110000110110;
#1 $display("%b", po);
# 1  pi=24'b100110000010001110100011;
#1 $display("%b", po);
# 1  pi=24'b100100100000101111011000;
#1 $display("%b", po);
# 1  pi=24'b110000000010010101110000;
#1 $display("%b", po);
# 1  pi=24'b111010011101000001111111;
#1 $display("%b", po);
# 1  pi=24'b011111110111000011001010;
#1 $display("%b", po);
# 1  pi=24'b000101000100100100011000;
#1 $display("%b", po);
# 1  pi=24'b011000001010001101100100;
#1 $display("%b", po);
# 1  pi=24'b011000110000001100010111;
#1 $display("%b", po);
# 1  pi=24'b101111100011000111111110;
#1 $display("%b", po);
# 1  pi=24'b010101010000000101111110;
#1 $display("%b", po);
# 1  pi=24'b011011010001000111011011;
#1 $display("%b", po);
# 1  pi=24'b010011010111111011011101;
#1 $display("%b", po);
# 1  pi=24'b000100010111101110001010;
#1 $display("%b", po);
# 1  pi=24'b111000101001001010011010;
#1 $display("%b", po);
# 1  pi=24'b101110001000000001010100;
#1 $display("%b", po);
# 1  pi=24'b000000010001010111110100;
#1 $display("%b", po);
# 1  pi=24'b110011100101011010010110;
#1 $display("%b", po);
# 1  pi=24'b000011100101110001101101;
#1 $display("%b", po);
# 1  pi=24'b010101001110001000111010;
#1 $display("%b", po);
# 1  pi=24'b001100111101000110100001;
#1 $display("%b", po);
# 1  pi=24'b001100010010111000001001;
#1 $display("%b", po);
# 1  pi=24'b111000000001100000010101;
#1 $display("%b", po);
# 1  pi=24'b110101100111101111110100;
#1 $display("%b", po);
# 1  pi=24'b010010111010011111100001;
#1 $display("%b", po);
# 1  pi=24'b011001011000100001110011;
#1 $display("%b", po);
# 1  pi=24'b000001110101100101111111;
#1 $display("%b", po);
# 1  pi=24'b101111111101111100110101;
#1 $display("%b", po);
# 1  pi=24'b001101000111000111110101;
#1 $display("%b", po);
# 1  pi=24'b101100101010110110001111;
#1 $display("%b", po);
# 1  pi=24'b001110110111000000010111;
#1 $display("%b", po);
# 1  pi=24'b101000011010100001001100;
#1 $display("%b", po);
# 1  pi=24'b101101111001110011011110;
#1 $display("%b", po);
# 1  pi=24'b011110011100100110101001;
#1 $display("%b", po);
# 1  pi=24'b101101001110001100000010;
#1 $display("%b", po);
# 1  pi=24'b001010011111111000011110;
#1 $display("%b", po);
# 1  pi=24'b110010000000000111001010;
#1 $display("%b", po);
# 1  pi=24'b110100000110100010101011;
#1 $display("%b", po);
# 1  pi=24'b111111111111010100011110;
#1 $display("%b", po);
# 1  pi=24'b000001100000011010100110;
#1 $display("%b", po);
# 1  pi=24'b011011100110110000000010;
#1 $display("%b", po);
# 1  pi=24'b011111010000111111101010;
#1 $display("%b", po);
# 1  pi=24'b000110001101000110100100;
#1 $display("%b", po);
# 1  pi=24'b010010110001100110000000;
#1 $display("%b", po);
# 1  pi=24'b111000001001000100000111;
#1 $display("%b", po);
# 1  pi=24'b011000101001101110000001;
#1 $display("%b", po);
# 1  pi=24'b001000111101101110001010;
#1 $display("%b", po);
# 1  pi=24'b101000101100100000010110;
#1 $display("%b", po);
# 1  pi=24'b010101000100101011000011;
#1 $display("%b", po);
# 1  pi=24'b010000011001001011100011;
#1 $display("%b", po);
# 1  pi=24'b011110101000111010100101;
#1 $display("%b", po);
# 1  pi=24'b000000011100100010111101;
#1 $display("%b", po);
# 1  pi=24'b111110011000111110110101;
#1 $display("%b", po);
# 1  pi=24'b010110110011100010110010;
#1 $display("%b", po);
# 1  pi=24'b011100000111101000110010;
#1 $display("%b", po);
# 1  pi=24'b111001011110011001000110;
#1 $display("%b", po);
# 1  pi=24'b011001001100111100111101;
#1 $display("%b", po);
# 1  pi=24'b010011111111000000111111;
#1 $display("%b", po);
# 1  pi=24'b000011000110111011110111;
#1 $display("%b", po);
# 1  pi=24'b110010010010010011100110;
#1 $display("%b", po);
# 1  pi=24'b001100011111000111100001;
#1 $display("%b", po);
# 1  pi=24'b110101100001001001110011;
#1 $display("%b", po);
# 1  pi=24'b100010101000111010000111;
#1 $display("%b", po);
# 1  pi=24'b110110000011101011101110;
#1 $display("%b", po);
# 1  pi=24'b001000001001010110000010;
#1 $display("%b", po);
# 1  pi=24'b101000100000001110100100;
#1 $display("%b", po);
# 1  pi=24'b001101111101000101000111;
#1 $display("%b", po);
# 1  pi=24'b000000100000110101110010;
#1 $display("%b", po);
# 1  pi=24'b101000111111101010000001;
#1 $display("%b", po);
# 1  pi=24'b110011011011011110001111;
#1 $display("%b", po);
# 1  pi=24'b101111000111100010111111;
#1 $display("%b", po);
# 1  pi=24'b000101101001101101001111;
#1 $display("%b", po);
# 1  pi=24'b000110011110101100111110;
#1 $display("%b", po);
# 1  pi=24'b010010010011010110110010;
#1 $display("%b", po);
# 1  pi=24'b000001000101110100100010;
#1 $display("%b", po);
# 1  pi=24'b100011101100110000111110;
#1 $display("%b", po);
# 1  pi=24'b010110000110011101101100;
#1 $display("%b", po);
# 1  pi=24'b001001100110101111111101;
#1 $display("%b", po);
# 1  pi=24'b001110001100001110110111;
#1 $display("%b", po);
# 1  pi=24'b010001011011001100100110;
#1 $display("%b", po);
# 1  pi=24'b001001011100011010101000;
#1 $display("%b", po);
# 1  pi=24'b011001101000111110010011;
#1 $display("%b", po);
# 1  pi=24'b001101011110000110011001;
#1 $display("%b", po);
# 1  pi=24'b001101100100101001001010;
#1 $display("%b", po);
# 1  pi=24'b010111000011000011000001;
#1 $display("%b", po);
# 1  pi=24'b100110100010111011110011;
#1 $display("%b", po);
# 1  pi=24'b110101010110111010001001;
#1 $display("%b", po);
# 1  pi=24'b010001111000011110001010;
#1 $display("%b", po);
# 1  pi=24'b001000101110110010101101;
#1 $display("%b", po);
# 1  pi=24'b010000010010110001110010;
#1 $display("%b", po);
# 1  pi=24'b001100111111001011001010;
#1 $display("%b", po);
# 1  pi=24'b000001110010001010011100;
#1 $display("%b", po);
# 1  pi=24'b011001110111000010110001;
#1 $display("%b", po);
# 1  pi=24'b010000111111000000011001;
#1 $display("%b", po);
# 1  pi=24'b111100110111110101101000;
#1 $display("%b", po);
# 1  pi=24'b000111011000110111011010;
#1 $display("%b", po);
# 1  pi=24'b010101000110001000011100;
#1 $display("%b", po);
# 1  pi=24'b100101001110101100100000;
#1 $display("%b", po);
# 1  pi=24'b000011111100011110110010;
#1 $display("%b", po);
# 1  pi=24'b010000101110001101110011;
#1 $display("%b", po);
# 1  pi=24'b100111111100001011010001;
#1 $display("%b", po);
# 1  pi=24'b000011010101001101010100;
#1 $display("%b", po);
# 1  pi=24'b010100001101111000000101;
#1 $display("%b", po);
# 1  pi=24'b001010001010110011011100;
#1 $display("%b", po);
# 1  pi=24'b111001010111001000111100;
#1 $display("%b", po);
# 1  pi=24'b111111100111100101110001;
#1 $display("%b", po);
# 1  pi=24'b111001111111001001111000;
#1 $display("%b", po);
# 1  pi=24'b000100000010000011111100;
#1 $display("%b", po);
# 1  pi=24'b100011010111010110011010;
#1 $display("%b", po);
# 1  pi=24'b011001101010110111100010;
#1 $display("%b", po);
# 1  pi=24'b001111001000110000010010;
#1 $display("%b", po);
# 1  pi=24'b000000101111000101110110;
#1 $display("%b", po);
# 1  pi=24'b101111101110001101000110;
#1 $display("%b", po);
# 1  pi=24'b110001010011110000000000;
#1 $display("%b", po);
# 1  pi=24'b111001111100000101101001;
#1 $display("%b", po);
# 1  pi=24'b100000111111010000111011;
#1 $display("%b", po);
# 1  pi=24'b100100000011100111011011;
#1 $display("%b", po);
# 1  pi=24'b001000101110101010011010;
#1 $display("%b", po);
# 1  pi=24'b100110101001110101000111;
#1 $display("%b", po);
# 1  pi=24'b000111101000101111011001;
#1 $display("%b", po);
# 1  pi=24'b101100010111000110011010;
#1 $display("%b", po);
# 1  pi=24'b110110100101000110110111;
#1 $display("%b", po);
# 1  pi=24'b110110101111001101110000;
#1 $display("%b", po);
# 1  pi=24'b010100101101000100110101;
#1 $display("%b", po);
# 1  pi=24'b111101110001001101101000;
#1 $display("%b", po);
# 1  pi=24'b101100110011100100110001;
#1 $display("%b", po);
# 1  pi=24'b100110111000000110101100;
#1 $display("%b", po);
# 1  pi=24'b111110000100001010111101;
#1 $display("%b", po);
# 1  pi=24'b011010110101100010011001;
#1 $display("%b", po);
# 1  pi=24'b100011010111001110110000;
#1 $display("%b", po);
# 1  pi=24'b001000000110011110100010;
#1 $display("%b", po);
# 1  pi=24'b011101001101000000101011;
#1 $display("%b", po);
# 1  pi=24'b110001000111001100011000;
#1 $display("%b", po);
# 1  pi=24'b101001001010000011011110;
#1 $display("%b", po);
# 1  pi=24'b101100100011000100111101;
#1 $display("%b", po);
# 1  pi=24'b001001011001110011000111;
#1 $display("%b", po);
# 1  pi=24'b001101111100100010111011;
#1 $display("%b", po);
# 1  pi=24'b001011100100010101110111;
#1 $display("%b", po);
# 1  pi=24'b110100101100100011000011;
#1 $display("%b", po);
# 1  pi=24'b101000001101011001000100;
#1 $display("%b", po);
# 1  pi=24'b101110010101100000100101;
#1 $display("%b", po);
# 1  pi=24'b100100001101100000101011;
#1 $display("%b", po);
# 1  pi=24'b000001001100011110110111;
#1 $display("%b", po);
# 1  pi=24'b100011101101111111101101;
#1 $display("%b", po);
# 1  pi=24'b101000000010001011110011;
#1 $display("%b", po);
# 1  pi=24'b011110101010000110010101;
#1 $display("%b", po);
# 1  pi=24'b001101101011100011011110;
#1 $display("%b", po);
# 1  pi=24'b110001111010000011101011;
#1 $display("%b", po);
# 1  pi=24'b000001010001111000011011;
#1 $display("%b", po);
# 1  pi=24'b001010001010000111010001;
#1 $display("%b", po);
# 1  pi=24'b101101010101111010100010;
#1 $display("%b", po);
# 1  pi=24'b100110101101100010110000;
#1 $display("%b", po);
# 1  pi=24'b000001100101111110110010;
#1 $display("%b", po);
# 1  pi=24'b101000101010010000010101;
#1 $display("%b", po);
# 1  pi=24'b000101010011011100111011;
#1 $display("%b", po);
# 1  pi=24'b101101110111101110011000;
#1 $display("%b", po);
# 1  pi=24'b000101001111110010010100;
#1 $display("%b", po);
# 1  pi=24'b010110110001111100100000;
#1 $display("%b", po);
# 1  pi=24'b000100011010101110110010;
#1 $display("%b", po);
# 1  pi=24'b010000000110001100000001;
#1 $display("%b", po);
# 1  pi=24'b011000001000111100010111;
#1 $display("%b", po);
# 1  pi=24'b011111011110011101010010;
#1 $display("%b", po);
# 1  pi=24'b011100010000110110010010;
#1 $display("%b", po);
# 1  pi=24'b100000100111011101011111;
#1 $display("%b", po);
# 1  pi=24'b011100010111100110101110;
#1 $display("%b", po);
# 1  pi=24'b000011110100111010100001;
#1 $display("%b", po);
# 1  pi=24'b011101100000110100001111;
#1 $display("%b", po);
# 1  pi=24'b100101111001101010011011;
#1 $display("%b", po);
# 1  pi=24'b000001000011111110111110;
#1 $display("%b", po);
# 1  pi=24'b110011001110100001010011;
#1 $display("%b", po);
# 1  pi=24'b000111000101010001100010;
#1 $display("%b", po);
# 1  pi=24'b001110110011011011010011;
#1 $display("%b", po);
# 1  pi=24'b011110000100010000111011;
#1 $display("%b", po);
# 1  pi=24'b010010001100011000000000;
#1 $display("%b", po);
# 1  pi=24'b011100101010110100111000;
#1 $display("%b", po);
# 1  pi=24'b011110111111011010101001;
#1 $display("%b", po);
# 1  pi=24'b010000011011000100101010;
#1 $display("%b", po);
# 1  pi=24'b011100111110010101100011;
#1 $display("%b", po);
# 1  pi=24'b111110000100101111110111;
#1 $display("%b", po);
# 1  pi=24'b011010000111101001001011;
#1 $display("%b", po);
# 1  pi=24'b111110111010011111110001;
#1 $display("%b", po);
# 1  pi=24'b110010110000110000000000;
#1 $display("%b", po);
# 1  pi=24'b100011101001000110101110;
#1 $display("%b", po);
# 1  pi=24'b000001000101110110001001;
#1 $display("%b", po);
# 1  pi=24'b001111101100110111011011;
#1 $display("%b", po);
# 1  pi=24'b010110101100001011100000;
#1 $display("%b", po);
# 1  pi=24'b001101011010010100111110;
#1 $display("%b", po);
# 1  pi=24'b000000000101000101010010;
#1 $display("%b", po);
# 1  pi=24'b010011110100100000100100;
#1 $display("%b", po);
# 1  pi=24'b111100101101000001010110;
#1 $display("%b", po);
# 1  pi=24'b010010000000111000011101;
#1 $display("%b", po);
# 1  pi=24'b110000010100111011000010;
#1 $display("%b", po);
# 1  pi=24'b110101001001110000101011;
#1 $display("%b", po);
# 1  pi=24'b000101011110010110000101;
#1 $display("%b", po);
# 1  pi=24'b101000001011000110100111;
#1 $display("%b", po);
# 1  pi=24'b100011110100001111100100;
#1 $display("%b", po);
# 1  pi=24'b110110010001001111100011;
#1 $display("%b", po);
# 1  pi=24'b011101110111011100111010;
#1 $display("%b", po);
# 1  pi=24'b010111111100100001011100;
#1 $display("%b", po);
# 1  pi=24'b111010110101001011010010;
#1 $display("%b", po);
# 1  pi=24'b110100011111111100011110;
#1 $display("%b", po);
# 1  pi=24'b000101101111000101100000;
#1 $display("%b", po);
# 1  pi=24'b011110000110111111010101;
#1 $display("%b", po);
# 1  pi=24'b111100101001101101110101;
#1 $display("%b", po);
# 1  pi=24'b110000110101111000100110;
#1 $display("%b", po);
# 1  pi=24'b001000011010101001101100;
#1 $display("%b", po);
# 1  pi=24'b011110100010011011101000;
#1 $display("%b", po);
# 1  pi=24'b010110101000000110011010;
#1 $display("%b", po);
# 1  pi=24'b110100111010110111111111;
#1 $display("%b", po);
# 1  pi=24'b010111000011100010000111;
#1 $display("%b", po);
# 1  pi=24'b101100011110010101111000;
#1 $display("%b", po);
# 1  pi=24'b110000000011111000011010;
#1 $display("%b", po);
# 1  pi=24'b010111001011101011100011;
#1 $display("%b", po);
# 1  pi=24'b000111111101111000100010;
#1 $display("%b", po);
# 1  pi=24'b011110000000100010111001;
#1 $display("%b", po);
# 1  pi=24'b001011011000000101111110;
#1 $display("%b", po);
# 1  pi=24'b111001000100011101011111;
#1 $display("%b", po);
# 1  pi=24'b111000011100111000111000;
#1 $display("%b", po);
# 1  pi=24'b010000110110110010000100;
#1 $display("%b", po);
# 1  pi=24'b000110101100000000010110;
#1 $display("%b", po);
# 1  pi=24'b101000110010000001101001;
#1 $display("%b", po);
# 1  pi=24'b000010101110101111100010;
#1 $display("%b", po);
# 1  pi=24'b010000100011100111111110;
#1 $display("%b", po);
# 1  pi=24'b100111110100110101110100;
#1 $display("%b", po);
# 1  pi=24'b000101000010110010111001;
#1 $display("%b", po);
# 1  pi=24'b111111011101011001100111;
#1 $display("%b", po);
# 1  pi=24'b001101001111101011001011;
#1 $display("%b", po);
# 1  pi=24'b100101000101000000111101;
#1 $display("%b", po);
# 1  pi=24'b111101001000100101110111;
#1 $display("%b", po);
# 1  pi=24'b001001100011111001111001;
#1 $display("%b", po);
# 1  pi=24'b110111011001001001100011;
#1 $display("%b", po);
# 1  pi=24'b011011101101100101100111;
#1 $display("%b", po);
# 1  pi=24'b110010000110001000011100;
#1 $display("%b", po);
# 1  pi=24'b001111100110001110101000;
#1 $display("%b", po);
# 1  pi=24'b110010101010011100101000;
#1 $display("%b", po);
# 1  pi=24'b101001111100100110001110;
#1 $display("%b", po);
# 1  pi=24'b100000011110001011010100;
#1 $display("%b", po);
# 1  pi=24'b011011010101111100011010;
#1 $display("%b", po);
# 1  pi=24'b110111010101011110110100;
#1 $display("%b", po);
# 1  pi=24'b000111001010010010011010;
#1 $display("%b", po);
# 1  pi=24'b111111001001110000011000;
#1 $display("%b", po);
# 1  pi=24'b100000100001010101000011;
#1 $display("%b", po);
# 1  pi=24'b111011111101111011000101;
#1 $display("%b", po);
# 1  pi=24'b011110101101011111011111;
#1 $display("%b", po);
# 1  pi=24'b101010010010110110111100;
#1 $display("%b", po);
# 1  pi=24'b000101001000111111110001;
#1 $display("%b", po);
# 1  pi=24'b101110110100011010110100;
#1 $display("%b", po);
# 1  pi=24'b110010010001001100111010;
#1 $display("%b", po);
# 1  pi=24'b000000010100110110000000;
#1 $display("%b", po);
# 1  pi=24'b111001111110100000101010;
#1 $display("%b", po);
# 1  pi=24'b001011010101011101111011;
#1 $display("%b", po);
# 1  pi=24'b010001000101010100010100;
#1 $display("%b", po);
# 1  pi=24'b110101000011001101011010;
#1 $display("%b", po);
# 1  pi=24'b011010011110000100010111;
#1 $display("%b", po);
# 1  pi=24'b010100001000000001001110;
#1 $display("%b", po);
# 1  pi=24'b111000110000001001101111;
#1 $display("%b", po);
# 1  pi=24'b101011001101111110110111;
#1 $display("%b", po);
# 1  pi=24'b001011100011001111010110;
#1 $display("%b", po);
# 1  pi=24'b100100001011010010000000;
#1 $display("%b", po);
# 1  pi=24'b010000001001011011011000;
#1 $display("%b", po);
# 1  pi=24'b010101101100010011010110;
#1 $display("%b", po);
# 1  pi=24'b110111010011100101011111;
#1 $display("%b", po);
# 1  pi=24'b111101101000010101100010;
#1 $display("%b", po);
# 1  pi=24'b100011011011000010010111;
#1 $display("%b", po);
# 1  pi=24'b101110001010101011000111;
#1 $display("%b", po);
# 1  pi=24'b111110000100000000100010;
#1 $display("%b", po);
# 1  pi=24'b111111001011101011111100;
#1 $display("%b", po);
# 1  pi=24'b000010011000101010100100;
#1 $display("%b", po);
# 1  pi=24'b010001110001101110001010;
#1 $display("%b", po);
# 1  pi=24'b010000101100100011010100;
#1 $display("%b", po);
# 1  pi=24'b100011010111111100010100;
#1 $display("%b", po);
# 1  pi=24'b110110101001001011101001;
#1 $display("%b", po);
# 1  pi=24'b111110011111100101110100;
#1 $display("%b", po);
# 1  pi=24'b001110110001000000000011;
#1 $display("%b", po);
# 1  pi=24'b001001110010011001100100;
#1 $display("%b", po);
# 1  pi=24'b111101011011101011010101;
#1 $display("%b", po);
# 1  pi=24'b100011110000001001001111;
#1 $display("%b", po);
# 1  pi=24'b010011100100111000001110;
#1 $display("%b", po);
# 1  pi=24'b111100000111000101110100;
#1 $display("%b", po);
# 1  pi=24'b110101111010100010110100;
#1 $display("%b", po);
# 1  pi=24'b011001011110001000101000;
#1 $display("%b", po);
# 1  pi=24'b100100101000110011101110;
#1 $display("%b", po);
# 1  pi=24'b000100110010011101110000;
#1 $display("%b", po);
# 1  pi=24'b011111101000010001001110;
#1 $display("%b", po);
# 1  pi=24'b001110100110000110010000;
#1 $display("%b", po);
# 1  pi=24'b111101101011101111011001;
#1 $display("%b", po);
# 1  pi=24'b110000010110111011100100;
#1 $display("%b", po);
# 1  pi=24'b011100111110110111010100;
#1 $display("%b", po);
# 1  pi=24'b100101001010010111001111;
#1 $display("%b", po);
# 1  pi=24'b000111010111100001100000;
#1 $display("%b", po);
# 1  pi=24'b110010100001110110111001;
#1 $display("%b", po);
# 1  pi=24'b011001100001001111111011;
#1 $display("%b", po);
# 1  pi=24'b100111000101000100110001;
#1 $display("%b", po);
# 1  pi=24'b110011110110101000010111;
#1 $display("%b", po);
# 1  pi=24'b010100101101011100110010;
#1 $display("%b", po);
# 1  pi=24'b000000101001100001001101;
#1 $display("%b", po);
# 1  pi=24'b001010001110101000101001;
#1 $display("%b", po);
# 1  pi=24'b111010110111000101101001;
#1 $display("%b", po);
# 1  pi=24'b000001000100010000000101;
#1 $display("%b", po);
# 1  pi=24'b100110100100011000110000;
#1 $display("%b", po);
# 1  pi=24'b100010100101111011000010;
#1 $display("%b", po);
# 1  pi=24'b000110101101010101101010;
#1 $display("%b", po);
# 1  pi=24'b101101111011110011011111;
#1 $display("%b", po);
# 1  pi=24'b000110110101000101000011;
#1 $display("%b", po);
# 1  pi=24'b010110101101010111100011;
#1 $display("%b", po);
# 1  pi=24'b101010000110100101011010;
#1 $display("%b", po);
# 1  pi=24'b110001011101101110110000;
#1 $display("%b", po);
# 1  pi=24'b000010010010111111111001;
#1 $display("%b", po);
# 1  pi=24'b010100111101011101011101;
#1 $display("%b", po);
# 1  pi=24'b111101000100011011001110;
#1 $display("%b", po);
# 1  pi=24'b010110011011001111000101;
#1 $display("%b", po);
# 1  pi=24'b000001110110010010010001;
#1 $display("%b", po);
# 1  pi=24'b011000101010100111011111;
#1 $display("%b", po);
# 1  pi=24'b001010110100101100000000;
#1 $display("%b", po);
# 1  pi=24'b101100101000000011101001;
#1 $display("%b", po);
# 1  pi=24'b011010100000011000001110;
#1 $display("%b", po);
# 1  pi=24'b010000100011100101011111;
#1 $display("%b", po);
# 1  pi=24'b000111111110011111110111;
#1 $display("%b", po);
# 1  pi=24'b000101101111101000111110;
#1 $display("%b", po);
# 1  pi=24'b011010000010011111010010;
#1 $display("%b", po);
# 1  pi=24'b010010000100010011011001;
#1 $display("%b", po);
# 1  pi=24'b001011110110110110111011;
#1 $display("%b", po);
# 1  pi=24'b001001000000100011101010;
#1 $display("%b", po);
# 1  pi=24'b111000000011111110000111;
#1 $display("%b", po);
# 1  pi=24'b110010000101010101101010;
#1 $display("%b", po);
# 1  pi=24'b011000011010110001010001;
#1 $display("%b", po);
# 1  pi=24'b101101111001001100100111;
#1 $display("%b", po);
# 1  pi=24'b101101010011001011111101;
#1 $display("%b", po);
# 1  pi=24'b111001011111010110111011;
#1 $display("%b", po);
# 1  pi=24'b100100101100111010011100;
#1 $display("%b", po);
# 1  pi=24'b101010100110110011011010;
#1 $display("%b", po);
# 1  pi=24'b100101101011010111110000;
#1 $display("%b", po);
# 1  pi=24'b001110011110110001011101;
#1 $display("%b", po);
# 1  pi=24'b011000010100000100001101;
#1 $display("%b", po);
# 1  pi=24'b100101011100101000100100;
#1 $display("%b", po);
# 1  pi=24'b001110010000000100110011;
#1 $display("%b", po);
# 1  pi=24'b011110110101110010110110;
#1 $display("%b", po);
# 1  pi=24'b011100111100010110000010;
#1 $display("%b", po);
# 1  pi=24'b110101010000101111000111;
#1 $display("%b", po);
# 1  pi=24'b001100001110100001000001;
#1 $display("%b", po);
# 1  pi=24'b100111010111100100101101;
#1 $display("%b", po);
# 1  pi=24'b011100100111110100000111;
#1 $display("%b", po);
# 1  pi=24'b100011111101111101001010;
#1 $display("%b", po);
# 1  pi=24'b101110010111100101001001;
#1 $display("%b", po);
# 1  pi=24'b010100000111011000110011;
#1 $display("%b", po);
# 1  pi=24'b011111000011000100101000;
#1 $display("%b", po);
# 1  pi=24'b111000000000011101001110;
#1 $display("%b", po);
# 1  pi=24'b011001001011101001100011;
#1 $display("%b", po);
# 1  pi=24'b110001011011000101001000;
#1 $display("%b", po);
# 1  pi=24'b001001001000010100110111;
#1 $display("%b", po);
# 1  pi=24'b101101101110010001101101;
#1 $display("%b", po);
# 1  pi=24'b000011110001100111101111;
#1 $display("%b", po);
# 1  pi=24'b111100011110101001011001;
#1 $display("%b", po);
# 1  pi=24'b110100111000110010100001;
#1 $display("%b", po);
# 1  pi=24'b111101001101111010111001;
#1 $display("%b", po);
# 1  pi=24'b100100010001001010101001;
#1 $display("%b", po);
# 1  pi=24'b101111001101100000110101;
#1 $display("%b", po);
# 1  pi=24'b011001001111010110111101;
#1 $display("%b", po);
# 1  pi=24'b010101110000000010110111;
#1 $display("%b", po);
# 1  pi=24'b110000110111101001101001;
#1 $display("%b", po);
# 1  pi=24'b111010000101011100000111;
#1 $display("%b", po);
# 1  pi=24'b100111001010100111110011;
#1 $display("%b", po);
# 1  pi=24'b010010110110101010110011;
#1 $display("%b", po);
# 1  pi=24'b011000101000000001010101;
#1 $display("%b", po);
# 1  pi=24'b000001011101011110001101;
#1 $display("%b", po);
# 1  pi=24'b000101110010000011010111;
#1 $display("%b", po);
# 1  pi=24'b110000111000011111001011;
#1 $display("%b", po);
# 1  pi=24'b011110011101101001001001;
#1 $display("%b", po);
# 1  pi=24'b001000011001101111011010;
#1 $display("%b", po);
# 1  pi=24'b001111010110011100010011;
#1 $display("%b", po);
# 1  pi=24'b000000111010000110100111;
#1 $display("%b", po);
# 1  pi=24'b000001000100000010000100;
#1 $display("%b", po);
# 1  pi=24'b010101001001011001010110;
#1 $display("%b", po);
# 1  pi=24'b100101110100000010100011;
#1 $display("%b", po);
# 1  pi=24'b010000010111001011000011;
#1 $display("%b", po);
# 1  pi=24'b110001001110000001010011;
#1 $display("%b", po);
# 1  pi=24'b010001101110101100010101;
#1 $display("%b", po);
# 1  pi=24'b100010011011100011000111;
#1 $display("%b", po);
# 1  pi=24'b001111001110000101001111;
#1 $display("%b", po);
# 1  pi=24'b100010111110010111000000;
#1 $display("%b", po);
# 1  pi=24'b110000110010111001110000;
#1 $display("%b", po);
# 1  pi=24'b111110100100010011000100;
#1 $display("%b", po);
# 1  pi=24'b000001000101101111101010;
#1 $display("%b", po);
# 1  pi=24'b111111110010111000011111;
#1 $display("%b", po);
# 1  pi=24'b111110101000100101000110;
#1 $display("%b", po);
# 1  pi=24'b011111011110101001111001;
#1 $display("%b", po);
# 1  pi=24'b011001010000001101110111;
#1 $display("%b", po);
# 1  pi=24'b100101110001100101111011;
#1 $display("%b", po);
# 1  pi=24'b010011000000000010011110;
#1 $display("%b", po);
# 1  pi=24'b110110100110101100000111;
#1 $display("%b", po);
# 1  pi=24'b011100011110000010011111;
#1 $display("%b", po);
# 1  pi=24'b111010001110010111111010;
#1 $display("%b", po);
# 1  pi=24'b100101000001100011001010;
#1 $display("%b", po);
# 1  pi=24'b001110101000000111010010;
#1 $display("%b", po);
# 1  pi=24'b111101001100011001010100;
#1 $display("%b", po);
# 1  pi=24'b110000000101110101111011;
#1 $display("%b", po);
# 1  pi=24'b101110100110000110000011;
#1 $display("%b", po);
# 1  pi=24'b101011010011001110011001;
#1 $display("%b", po);
# 1  pi=24'b101011101010011111010011;
#1 $display("%b", po);
# 1  pi=24'b000110011101001001001000;
#1 $display("%b", po);
# 1  pi=24'b101011000011010011001001;
#1 $display("%b", po);
# 1  pi=24'b100100001011001111001100;
#1 $display("%b", po);
# 1  pi=24'b100110001100100000000011;
#1 $display("%b", po);
# 1  pi=24'b000110100101111011000111;
#1 $display("%b", po);
# 1  pi=24'b000110101010100010111110;
#1 $display("%b", po);
# 1  pi=24'b000000100110010001011110;
#1 $display("%b", po);
# 1  pi=24'b100110101100110011011010;
#1 $display("%b", po);
# 1  pi=24'b000010111010011000001010;
#1 $display("%b", po);
# 1  pi=24'b111011111000100101001010;
#1 $display("%b", po);
# 1  pi=24'b010011011110100101010111;
#1 $display("%b", po);
# 1  pi=24'b000001110110100100011111;
#1 $display("%b", po);
# 1  pi=24'b000111100101110100000011;
#1 $display("%b", po);
# 1  pi=24'b001001101011010111101010;
#1 $display("%b", po);
# 1  pi=24'b010010000110000100100000;
#1 $display("%b", po);
# 1  pi=24'b000101011110001001010001;
#1 $display("%b", po);
# 1  pi=24'b100100101101010011100110;
#1 $display("%b", po);
# 1  pi=24'b011011110011000110110011;
#1 $display("%b", po);
# 1  pi=24'b010100011111001100110111;
#1 $display("%b", po);
# 1  pi=24'b110010001110001010001010;
#1 $display("%b", po);
# 1  pi=24'b000000111111010100111101;
#1 $display("%b", po);
# 1  pi=24'b101101011101000001011111;
#1 $display("%b", po);
# 1  pi=24'b100101110001100010110010;
#1 $display("%b", po);
# 1  pi=24'b101110011010001011000110;
#1 $display("%b", po);
# 1  pi=24'b011000000010100000111100;
#1 $display("%b", po);
# 1  pi=24'b001100001001000100011010;
#1 $display("%b", po);
# 1  pi=24'b101000101100101110010110;
#1 $display("%b", po);
# 1  pi=24'b100001110111110100001101;
#1 $display("%b", po);
# 1  pi=24'b010110001001010011111110;
#1 $display("%b", po);
# 1  pi=24'b101100010111101010101110;
#1 $display("%b", po);
# 1  pi=24'b010110100111001001110010;
#1 $display("%b", po);
# 1  pi=24'b100000010001010010100100;
#1 $display("%b", po);
# 1  pi=24'b100000101110100000110101;
#1 $display("%b", po);
# 1  pi=24'b001000101110010110110100;
#1 $display("%b", po);
# 1  pi=24'b100111111110101010001111;
#1 $display("%b", po);
# 1  pi=24'b011110010101011101011111;
#1 $display("%b", po);
# 1  pi=24'b100001111110011010111000;
#1 $display("%b", po);
# 1  pi=24'b110011011110110011011000;
#1 $display("%b", po);
# 1  pi=24'b000001101110100110001011;
#1 $display("%b", po);
# 1  pi=24'b011101001101100010001001;
#1 $display("%b", po);
# 1  pi=24'b101011110001011101110110;
#1 $display("%b", po);
# 1  pi=24'b000100111010010111111101;
#1 $display("%b", po);
# 1  pi=24'b101101011010111111011000;
#1 $display("%b", po);
# 1  pi=24'b000100000001001000010100;
#1 $display("%b", po);
# 1  pi=24'b011100000001111101111110;
#1 $display("%b", po);
# 1  pi=24'b001011010100110001011010;
#1 $display("%b", po);
# 1  pi=24'b001101011110010011011101;
#1 $display("%b", po);
# 1  pi=24'b101100111101101010011101;
#1 $display("%b", po);
# 1  pi=24'b110100111011011100000000;
#1 $display("%b", po);
# 1  pi=24'b010100011000011001111100;
#1 $display("%b", po);
# 1  pi=24'b101101101111001011000101;
#1 $display("%b", po);
# 1  pi=24'b011101110000011011011001;
#1 $display("%b", po);
# 1  pi=24'b000011010010011001110010;
#1 $display("%b", po);
# 1  pi=24'b011100010001010110011100;
#1 $display("%b", po);
# 1  pi=24'b100101101101101111010000;
#1 $display("%b", po);
# 1  pi=24'b000011011011110101110110;
#1 $display("%b", po);
# 1  pi=24'b101001110100100010010000;
#1 $display("%b", po);
# 1  pi=24'b101010000010110101100000;
#1 $display("%b", po);
# 1  pi=24'b010011100110000100010110;
#1 $display("%b", po);
# 1  pi=24'b111010011100000000111101;
#1 $display("%b", po);
# 1  pi=24'b100011110110010001101111;
#1 $display("%b", po);
# 1  pi=24'b011111010101000000011011;
#1 $display("%b", po);
# 1  pi=24'b110110010111001111111100;
#1 $display("%b", po);
# 1  pi=24'b000001110111101110100110;
#1 $display("%b", po);
# 1  pi=24'b010101000100101010101111;
#1 $display("%b", po);
# 1  pi=24'b011110010000000110110001;
#1 $display("%b", po);
# 1  pi=24'b011110111010011010101111;
#1 $display("%b", po);
# 1  pi=24'b011000111100000011110010;
#1 $display("%b", po);
# 1  pi=24'b000111001011011011111101;
#1 $display("%b", po);
# 1  pi=24'b000011010101111000101111;
#1 $display("%b", po);
# 1  pi=24'b101001100011011011001100;
#1 $display("%b", po);
# 1  pi=24'b000000001100101111101111;
#1 $display("%b", po);
# 1  pi=24'b010010011001101010111101;
#1 $display("%b", po);
# 1  pi=24'b100011100111101001000000;
#1 $display("%b", po);
# 1  pi=24'b010101010110110110010010;
#1 $display("%b", po);
# 1  pi=24'b000110100111110011100001;
#1 $display("%b", po);
# 1  pi=24'b010011100011011010001100;
#1 $display("%b", po);
# 1  pi=24'b101100101111101010101011;
#1 $display("%b", po);
# 1  pi=24'b000100100111000110010111;
#1 $display("%b", po);
# 1  pi=24'b000111011010100101110110;
#1 $display("%b", po);
# 1  pi=24'b110010000000011011110110;
#1 $display("%b", po);
# 1  pi=24'b110100011110110010011011;
#1 $display("%b", po);
# 1  pi=24'b010101101100000000111111;
#1 $display("%b", po);
# 1  pi=24'b110100100100011010101110;
#1 $display("%b", po);
# 1  pi=24'b011000100111110011111011;
#1 $display("%b", po);
# 1  pi=24'b110000001101100010101010;
#1 $display("%b", po);
# 1  pi=24'b011101110110000111101100;
#1 $display("%b", po);
# 1  pi=24'b101111011111100001010100;
#1 $display("%b", po);
# 1  pi=24'b000000110110001111011110;
#1 $display("%b", po);
# 1  pi=24'b011111100011110101111111;
#1 $display("%b", po);
# 1  pi=24'b011001110101111111001010;
#1 $display("%b", po);
# 1  pi=24'b101000010111000001110111;
#1 $display("%b", po);
# 1  pi=24'b101000101110101011000101;
#1 $display("%b", po);
# 1  pi=24'b000010110010111101011101;
#1 $display("%b", po);
# 1  pi=24'b010110001001011101110001;
#1 $display("%b", po);
# 1  pi=24'b000100110100010001101000;
#1 $display("%b", po);
# 1  pi=24'b010010101110110010110000;
#1 $display("%b", po);
# 1  pi=24'b110110010110010011011011;
#1 $display("%b", po);
# 1  pi=24'b100011011101101101001011;
#1 $display("%b", po);
# 1  pi=24'b000110101111011010001001;
#1 $display("%b", po);
# 1  pi=24'b000001101101101010111000;
#1 $display("%b", po);
# 1  pi=24'b010001100010110011110001;
#1 $display("%b", po);
# 1  pi=24'b001011010001101000111101;
#1 $display("%b", po);
# 1  pi=24'b111110110000001110101100;
#1 $display("%b", po);
# 1  pi=24'b010100100010110011111000;
#1 $display("%b", po);
# 1  pi=24'b111001111010010000111100;
#1 $display("%b", po);
# 1  pi=24'b101010001101001001101001;
#1 $display("%b", po);
# 1  pi=24'b010111111100001110111110;
#1 $display("%b", po);
# 1  pi=24'b101010100111101010110100;
#1 $display("%b", po);
# 1  pi=24'b010110010111100110110100;
#1 $display("%b", po);
# 1  pi=24'b011100011110110111011011;
#1 $display("%b", po);
# 1  pi=24'b010110111001000011111010;
#1 $display("%b", po);
# 1  pi=24'b000001001011010110011111;
#1 $display("%b", po);
# 1  pi=24'b010011001000010011100110;
#1 $display("%b", po);
# 1  pi=24'b100111110101001100011101;
#1 $display("%b", po);
# 1  pi=24'b000001011000110111011000;
#1 $display("%b", po);
# 1  pi=24'b100001111000000001010110;
#1 $display("%b", po);
# 1  pi=24'b111110000100101000110011;
#1 $display("%b", po);
# 1  pi=24'b111101101010001101110010;
#1 $display("%b", po);
# 1  pi=24'b010001111011000111100000;
#1 $display("%b", po);
# 1  pi=24'b101111011101101111000101;
#1 $display("%b", po);
# 1  pi=24'b011111000101000100110100;
#1 $display("%b", po);
# 1  pi=24'b110100110110001010100001;
#1 $display("%b", po);
# 1  pi=24'b000000100001110011110101;
#1 $display("%b", po);
# 1  pi=24'b110100011110001101001111;
#1 $display("%b", po);
# 1  pi=24'b110100101100111001111000;
#1 $display("%b", po);
# 1  pi=24'b111011101010111000111101;
#1 $display("%b", po);
# 1  pi=24'b001100001100001101011101;
#1 $display("%b", po);
# 1  pi=24'b101000011001111000101101;
#1 $display("%b", po);
# 1  pi=24'b110111111000100101011111;
#1 $display("%b", po);
# 1  pi=24'b111100010110101111011000;
#1 $display("%b", po);
# 1  pi=24'b110101000110010010100110;
#1 $display("%b", po);
# 1  pi=24'b110011011011000001100101;
#1 $display("%b", po);
# 1  pi=24'b100101000011000010111101;
#1 $display("%b", po);
# 1  pi=24'b001111001111010011011001;
#1 $display("%b", po);
# 1  pi=24'b100100011000001111001011;
#1 $display("%b", po);
# 1  pi=24'b101000101010010100001001;
#1 $display("%b", po);
# 1  pi=24'b100011001011101000010010;
#1 $display("%b", po);
# 1  pi=24'b000101111101010111010101;
#1 $display("%b", po);
# 1  pi=24'b101000011101101111010111;
#1 $display("%b", po);
# 1  pi=24'b100001000001111011011111;
#1 $display("%b", po);
# 1  pi=24'b010101100000100011110000;
#1 $display("%b", po);
# 1  pi=24'b110111011000110001101011;
#1 $display("%b", po);
# 1  pi=24'b110010101101011110010111;
#1 $display("%b", po);
# 1  pi=24'b001100101001001110011011;
#1 $display("%b", po);
# 1  pi=24'b100110111111000011010011;
#1 $display("%b", po);
# 1  pi=24'b100001110000101000011111;
#1 $display("%b", po);
# 1  pi=24'b011001000100101011011001;
#1 $display("%b", po);
# 1  pi=24'b111000000100111011111101;
#1 $display("%b", po);
# 1  pi=24'b000101110111101010111101;
#1 $display("%b", po);
# 1  pi=24'b100110000010110000100101;
#1 $display("%b", po);
# 1  pi=24'b001000011111001001100010;
#1 $display("%b", po);
# 1  pi=24'b111101010010110100011001;
#1 $display("%b", po);
# 1  pi=24'b101010100101000100011011;
#1 $display("%b", po);
# 1  pi=24'b000111001010010011011101;
#1 $display("%b", po);
# 1  pi=24'b100001110000100110101100;
#1 $display("%b", po);
# 1  pi=24'b111000010001111100110000;
#1 $display("%b", po);
# 1  pi=24'b011100101101010000101011;
#1 $display("%b", po);
# 1  pi=24'b001101111101010101110101;
#1 $display("%b", po);
# 1  pi=24'b110100001010010111101111;
#1 $display("%b", po);
# 1  pi=24'b011001100100000111110001;
#1 $display("%b", po);
# 1  pi=24'b000000000110100010101100;
#1 $display("%b", po);
# 1  pi=24'b110100001100010011010011;
#1 $display("%b", po);
# 1  pi=24'b010000010001001100100110;
#1 $display("%b", po);
# 1  pi=24'b100110101110100111000011;
#1 $display("%b", po);
# 1  pi=24'b011100001001000101100001;
#1 $display("%b", po);
# 1  pi=24'b010001010101101110011001;
#1 $display("%b", po);
# 1  pi=24'b010000101110000011101110;
#1 $display("%b", po);
# 1  pi=24'b101110001011011100111000;
#1 $display("%b", po);
# 1  pi=24'b010001100010000100010011;
#1 $display("%b", po);
# 1  pi=24'b000111000101110111111101;
#1 $display("%b", po);
# 1  pi=24'b000010100100101111110100;
#1 $display("%b", po);
# 1  pi=24'b010001001100101101000001;
#1 $display("%b", po);
# 1  pi=24'b011100001100000010010010;
#1 $display("%b", po);
# 1  pi=24'b011110010010010110110011;
#1 $display("%b", po);
# 1  pi=24'b110000000111000111011010;
#1 $display("%b", po);
# 1  pi=24'b000001011100111111011110;
#1 $display("%b", po);
# 1  pi=24'b101000111101101000010011;
#1 $display("%b", po);
# 1  pi=24'b100000110100100010110110;
#1 $display("%b", po);
# 1  pi=24'b110000000000111011111111;
#1 $display("%b", po);
# 1  pi=24'b011000101011000010111111;
#1 $display("%b", po);
# 1  pi=24'b111100101000000000100010;
#1 $display("%b", po);
# 1  pi=24'b010000011000110011000011;
#1 $display("%b", po);
# 1  pi=24'b010001111101011111110000;
#1 $display("%b", po);
# 1  pi=24'b110101111011010101100101;
#1 $display("%b", po);
# 1  pi=24'b000000011101010000010111;
#1 $display("%b", po);
# 1  pi=24'b111111110110010111000000;
#1 $display("%b", po);
# 1  pi=24'b011000000101111100101100;
#1 $display("%b", po);
# 1  pi=24'b100101011001000000001100;
#1 $display("%b", po);
# 1  pi=24'b010111011011010010010011;
#1 $display("%b", po);
# 1  pi=24'b000010000110100010100101;
#1 $display("%b", po);
# 1  pi=24'b101001100011101010000000;
#1 $display("%b", po);
# 1  pi=24'b110011000010100010101111;
#1 $display("%b", po);
# 1  pi=24'b000010010010011010110001;
#1 $display("%b", po);
# 1  pi=24'b101000001010011001110100;
#1 $display("%b", po);
# 1  pi=24'b110111011110101100110011;
#1 $display("%b", po);
# 1  pi=24'b110010101000111111110111;
#1 $display("%b", po);
# 1  pi=24'b011101011010001001001101;
#1 $display("%b", po);
# 1  pi=24'b110100101110000100000101;
#1 $display("%b", po);
# 1  pi=24'b110011110000010110100110;
#1 $display("%b", po);
# 1  pi=24'b100100100001110000011100;
#1 $display("%b", po);
# 1  pi=24'b111011101111010101001011;
#1 $display("%b", po);
# 1  pi=24'b111000011010000010001101;
#1 $display("%b", po);
# 1  pi=24'b101001100101101001101110;
#1 $display("%b", po);
# 1  pi=24'b100100011001100110010000;
#1 $display("%b", po);
# 1  pi=24'b101011111000001100001111;
#1 $display("%b", po);
# 1  pi=24'b010011110000011111010111;
#1 $display("%b", po);
# 1  pi=24'b010000011001101011010011;
#1 $display("%b", po);
# 1  pi=24'b001010110110010001100100;
#1 $display("%b", po);
# 1  pi=24'b100011100101101000000001;
#1 $display("%b", po);
# 1  pi=24'b111110101101110010001100;
#1 $display("%b", po);
# 1  pi=24'b001001011011100000100001;
#1 $display("%b", po);
# 1  pi=24'b001000010101001000101100;
#1 $display("%b", po);
# 1  pi=24'b101101101011111111010100;
#1 $display("%b", po);
# 1  pi=24'b010101000110010011100000;
#1 $display("%b", po);
# 1  pi=24'b000011110101101111011001;
#1 $display("%b", po);
# 1  pi=24'b010100010110110011001011;
#1 $display("%b", po);
# 1  pi=24'b011111110011010111010001;
#1 $display("%b", po);
# 1  pi=24'b111101100000010010001111;
#1 $display("%b", po);
# 1  pi=24'b110001110001111000001111;
#1 $display("%b", po);
# 1  pi=24'b110001010001100101000111;
#1 $display("%b", po);
# 1  pi=24'b111111100000100011111001;
#1 $display("%b", po);
# 1  pi=24'b011110011000101110111000;
#1 $display("%b", po);
# 1  pi=24'b100111110001000110010110;
#1 $display("%b", po);
# 1  pi=24'b001000010101110010101111;
#1 $display("%b", po);
# 1  pi=24'b000000011111010111010010;
#1 $display("%b", po);
# 1  pi=24'b101100010111101010101000;
#1 $display("%b", po);
# 1  pi=24'b110111110010111001110100;
#1 $display("%b", po);
# 1  pi=24'b111001111111000100110000;
#1 $display("%b", po);
# 1  pi=24'b001111110000101011010010;
#1 $display("%b", po);
# 1  pi=24'b101010010100100001010101;
#1 $display("%b", po);
# 1  pi=24'b000010000110001010011011;
#1 $display("%b", po);
# 1  pi=24'b100000101100110000000100;
#1 $display("%b", po);
# 1  pi=24'b001000110100000000110100;
#1 $display("%b", po);
# 1  pi=24'b100010101001010101100111;
#1 $display("%b", po);
# 1  pi=24'b101100010000110000111001;
#1 $display("%b", po);
# 1  pi=24'b000110110100111101100011;
#1 $display("%b", po);
# 1  pi=24'b101000110110011110100000;
#1 $display("%b", po);
# 1  pi=24'b010011010100010111100011;
#1 $display("%b", po);
# 1  pi=24'b011110001101111101010111;
#1 $display("%b", po);
# 1  pi=24'b011111101011100000101110;
#1 $display("%b", po);
# 1  pi=24'b110111100100100011001000;
#1 $display("%b", po);
# 1  pi=24'b100101010100111010100001;
#1 $display("%b", po);
# 1  pi=24'b110100000010100110011111;
#1 $display("%b", po);
# 1  pi=24'b010011110110101101100100;
#1 $display("%b", po);
# 1  pi=24'b000001100101011011100110;
#1 $display("%b", po);
# 1  pi=24'b111001111101001001110011;
#1 $display("%b", po);
# 1  pi=24'b110011011010010110101001;
#1 $display("%b", po);
# 1  pi=24'b111110010001101010010011;
#1 $display("%b", po);
# 1  pi=24'b111010000011100011100101;
#1 $display("%b", po);
# 1  pi=24'b010100011000101100110100;
#1 $display("%b", po);
# 1  pi=24'b001001110100100001010010;
#1 $display("%b", po);
# 1  pi=24'b001100000101101110011100;
#1 $display("%b", po);
# 1  pi=24'b110001011110001011100101;
#1 $display("%b", po);
# 1  pi=24'b000111111111100110100110;
#1 $display("%b", po);
# 1  pi=24'b111101001001110101011111;
#1 $display("%b", po);
# 1  pi=24'b101010100000111001111101;
#1 $display("%b", po);
# 1  pi=24'b011111010001100100010111;
#1 $display("%b", po);
# 1  pi=24'b001101100000100000101110;
#1 $display("%b", po);
# 1  pi=24'b000101100111000001001001;
#1 $display("%b", po);
# 1  pi=24'b111110110011101101101111;
#1 $display("%b", po);
# 1  pi=24'b101101111010111011010011;
#1 $display("%b", po);
# 1  pi=24'b010010011000101001001010;
#1 $display("%b", po);
# 1  pi=24'b101111000100111100111111;
#1 $display("%b", po);
# 1  pi=24'b101001000000000001110101;
#1 $display("%b", po);
# 1  pi=24'b010111100011100101001001;
#1 $display("%b", po);
# 1  pi=24'b111100110111110011110001;
#1 $display("%b", po);
# 1  pi=24'b100010111000001010001011;
#1 $display("%b", po);
# 1  pi=24'b001111101101100110110100;
#1 $display("%b", po);
# 1  pi=24'b011111110101111100111111;
#1 $display("%b", po);
# 1  pi=24'b110010111100010000110001;
#1 $display("%b", po);
# 1  pi=24'b100011100101001001101110;
#1 $display("%b", po);
# 1  pi=24'b111111000000010000000000;
#1 $display("%b", po);
# 1  pi=24'b001010101010100001100101;
#1 $display("%b", po);
# 1  pi=24'b000010010001001010000010;
#1 $display("%b", po);
# 1  pi=24'b011010101000100000000010;
#1 $display("%b", po);
# 1  pi=24'b001000000111000110100110;
#1 $display("%b", po);
# 1  pi=24'b011011001000100001111101;
#1 $display("%b", po);
# 1  pi=24'b010100001111100000100100;
#1 $display("%b", po);
# 1  pi=24'b110001101110011101010010;
#1 $display("%b", po);
# 1  pi=24'b110001000111000010010110;
#1 $display("%b", po);
# 1  pi=24'b110110011110000011111110;
#1 $display("%b", po);
# 1  pi=24'b010100101110101001000000;
#1 $display("%b", po);
# 1  pi=24'b100010100111001101011000;
#1 $display("%b", po);
# 1  pi=24'b011111010011100111100001;
#1 $display("%b", po);
# 1  pi=24'b110010011111010110111111;
#1 $display("%b", po);
# 1  pi=24'b010101001010001100100010;
#1 $display("%b", po);
# 1  pi=24'b001011001110000011010000;
#1 $display("%b", po);
# 1  pi=24'b101110101101001111111111;
#1 $display("%b", po);
# 1  pi=24'b100111111010011010110100;
#1 $display("%b", po);
# 1  pi=24'b010000000011010111101011;
#1 $display("%b", po);
# 1  pi=24'b000100110001011011001101;
#1 $display("%b", po);
# 1  pi=24'b001000100011000001110111;
#1 $display("%b", po);
# 1  pi=24'b000101110000110101111000;
#1 $display("%b", po);
# 1  pi=24'b010011011001010110110110;
#1 $display("%b", po);
# 1  pi=24'b100110100110000110101001;
#1 $display("%b", po);
# 1  pi=24'b001101011101000010110001;
#1 $display("%b", po);
# 1  pi=24'b100101100011000001111011;
#1 $display("%b", po);
# 1  pi=24'b111100010000111001110101;
#1 $display("%b", po);
# 1  pi=24'b100100101110111100101010;
#1 $display("%b", po);
# 1  pi=24'b001000110010111101000000;
#1 $display("%b", po);
# 1  pi=24'b010110001110101111001011;
#1 $display("%b", po);
# 1  pi=24'b101001000111000011010100;
#1 $display("%b", po);
# 1  pi=24'b110001110001011100110100;
#1 $display("%b", po);
# 1  pi=24'b000011001010111111100010;
#1 $display("%b", po);
# 1  pi=24'b101110100001000000011111;
#1 $display("%b", po);
# 1  pi=24'b111010010001110000001101;
#1 $display("%b", po);
# 1  pi=24'b100010101110101100000111;
#1 $display("%b", po);
# 1  pi=24'b101100101110111010111010;
#1 $display("%b", po);
# 1  pi=24'b010010011000101010100011;
#1 $display("%b", po);
# 1  pi=24'b010010000111000011100000;
#1 $display("%b", po);
# 1  pi=24'b010010111011011010111000;
#1 $display("%b", po);
# 1  pi=24'b111001010101110101111000;
#1 $display("%b", po);
# 1  pi=24'b101010101111101011111011;
#1 $display("%b", po);
# 1  pi=24'b111010000101100110010000;
#1 $display("%b", po);
# 1  pi=24'b000110100100101101000001;
#1 $display("%b", po);
# 1  pi=24'b101100010100001110001001;
#1 $display("%b", po);
# 1  pi=24'b010010001011001110111010;
#1 $display("%b", po);
# 1  pi=24'b011111001100010001001011;
#1 $display("%b", po);
# 1  pi=24'b100111100110010111001111;
#1 $display("%b", po);
# 1  pi=24'b101011100100011011111011;
#1 $display("%b", po);
# 1  pi=24'b111011011001011110110010;
#1 $display("%b", po);
# 1  pi=24'b101110101010011011100011;
#1 $display("%b", po);
# 1  pi=24'b100111101000111010001000;
#1 $display("%b", po);
# 1  pi=24'b111011011000100001010110;
#1 $display("%b", po);
# 1  pi=24'b011001101111010100000110;
#1 $display("%b", po);
# 1  pi=24'b001110101001010111010100;
#1 $display("%b", po);
# 1  pi=24'b111011001111110011100100;
#1 $display("%b", po);
# 1  pi=24'b010101010000000011101101;
#1 $display("%b", po);
# 1  pi=24'b100111011000101011011101;
#1 $display("%b", po);
# 1  pi=24'b011101110101111010000110;
#1 $display("%b", po);
# 1  pi=24'b000110111000000110010110;
#1 $display("%b", po);
# 1  pi=24'b100011000001110001000011;
#1 $display("%b", po);
# 1  pi=24'b010000110100111001100000;
#1 $display("%b", po);
# 1  pi=24'b010111111000011010011010;
#1 $display("%b", po);
# 1  pi=24'b111111010111110010100011;
#1 $display("%b", po);
# 1  pi=24'b101111011110101010101100;
#1 $display("%b", po);
# 1  pi=24'b101000010100011011111011;
#1 $display("%b", po);
# 1  pi=24'b101010011100101010110110;
#1 $display("%b", po);
# 1  pi=24'b101101100000101100010001;
#1 $display("%b", po);
# 1  pi=24'b110000011010001000011000;
#1 $display("%b", po);
# 1  pi=24'b011110001100010001110111;
#1 $display("%b", po);
# 1  pi=24'b101001101110100100101001;
#1 $display("%b", po);
# 1  pi=24'b000011011010101000110100;
#1 $display("%b", po);
# 1  pi=24'b000111010111011111011010;
#1 $display("%b", po);
# 1  pi=24'b001010110010010010010110;
#1 $display("%b", po);
# 1  pi=24'b100010110011010011111101;
#1 $display("%b", po);
# 1  pi=24'b110011010111000110100001;
#1 $display("%b", po);
# 1  pi=24'b110010111101101100010001;
#1 $display("%b", po);
# 1  pi=24'b111100011001100010011101;
#1 $display("%b", po);
# 1  pi=24'b011110001101011101100010;
#1 $display("%b", po);
# 1  pi=24'b010100000100110110111011;
#1 $display("%b", po);
# 1  pi=24'b001000110101101101010111;
#1 $display("%b", po);
# 1  pi=24'b011001010101000100110000;
#1 $display("%b", po);
# 1  pi=24'b011000010010001100011110;
#1 $display("%b", po);
# 1  pi=24'b110101011100000011100110;
#1 $display("%b", po);
# 1  pi=24'b110010010101100001111001;
#1 $display("%b", po);
# 1  pi=24'b010101111000100101001100;
#1 $display("%b", po);
# 1  pi=24'b010000001001111110111011;
#1 $display("%b", po);
# 1  pi=24'b011001110000100101110011;
#1 $display("%b", po);
# 1  pi=24'b111111100011011010001001;
#1 $display("%b", po);
# 1  pi=24'b110100010011010000010010;
#1 $display("%b", po);
# 1  pi=24'b110111010100111001011111;
#1 $display("%b", po);
# 1  pi=24'b110101100010101111100000;
#1 $display("%b", po);
# 1  pi=24'b010000000101101000111100;
#1 $display("%b", po);
# 1  pi=24'b110111001011000110111100;
#1 $display("%b", po);
# 1  pi=24'b011010111100000011110001;
#1 $display("%b", po);
# 1  pi=24'b010101100000111101011101;
#1 $display("%b", po);
# 1  pi=24'b111111011111100011110100;
#1 $display("%b", po);
# 1  pi=24'b011101010000001001000011;
#1 $display("%b", po);
# 1  pi=24'b100101110111011100100000;
#1 $display("%b", po);
# 1  pi=24'b111101100100111110111001;
#1 $display("%b", po);
# 1  pi=24'b111000001010000010000111;
#1 $display("%b", po);
# 1  pi=24'b011100110011001110111111;
#1 $display("%b", po);
# 1  pi=24'b000000100101011111100111;
#1 $display("%b", po);
# 1  pi=24'b010011011000101010001010;
#1 $display("%b", po);
# 1  pi=24'b000111100000001010000001;
#1 $display("%b", po);
# 1  pi=24'b000100011010111011010100;
#1 $display("%b", po);
# 1  pi=24'b000101100011100011000011;
#1 $display("%b", po);
# 1  pi=24'b001011001100011111111100;
#1 $display("%b", po);
# 1  pi=24'b101000101111100001010000;
#1 $display("%b", po);
# 1  pi=24'b001010000001010010001011;
#1 $display("%b", po);
# 1  pi=24'b010101101101001000001100;
#1 $display("%b", po);
# 1  pi=24'b000001101100110001000000;
#1 $display("%b", po);
# 1  pi=24'b111100001101011100100110;
#1 $display("%b", po);
# 1  pi=24'b001000011110011011011011;
#1 $display("%b", po);
# 1  pi=24'b000101000001001001001100;
#1 $display("%b", po);
# 1  pi=24'b010100001010111011010001;
#1 $display("%b", po);
# 1  pi=24'b000100010100001011011000;
#1 $display("%b", po);
# 1  pi=24'b101000001000011101101011;
#1 $display("%b", po);
# 1  pi=24'b001000001010111001000110;
#1 $display("%b", po);
# 1  pi=24'b111101100011100111001101;
#1 $display("%b", po);
# 1  pi=24'b101101100100001010010000;
#1 $display("%b", po);
# 1  pi=24'b100100111111001110100000;
#1 $display("%b", po);
# 1  pi=24'b111100111000100001100010;
#1 $display("%b", po);
# 1  pi=24'b010010011010101000010010;
#1 $display("%b", po);
# 1  pi=24'b000010101111101000011110;
#1 $display("%b", po);
# 1  pi=24'b010111100111000100001111;
#1 $display("%b", po);
# 1  pi=24'b001111010001011111110110;
#1 $display("%b", po);
# 1  pi=24'b011001101001101100011100;
#1 $display("%b", po);
# 1  pi=24'b111110110010111011001110;
#1 $display("%b", po);
# 1  pi=24'b111101000011100010110001;
#1 $display("%b", po);
# 1  pi=24'b100001101111100101010000;
#1 $display("%b", po);
# 1  pi=24'b100001011000011010011100;
#1 $display("%b", po);
# 1  pi=24'b010111101110001100000100;
#1 $display("%b", po);
# 1  pi=24'b000101111111010110000010;
#1 $display("%b", po);
# 1  pi=24'b110100100011000100110000;
#1 $display("%b", po);
# 1  pi=24'b000111110101000111100001;
#1 $display("%b", po);
# 1  pi=24'b000101110010101101010011;
#1 $display("%b", po);
# 1  pi=24'b100101100001011111000101;
#1 $display("%b", po);
# 1  pi=24'b010010001010011000001101;
#1 $display("%b", po);
# 1  pi=24'b011000010100011110011010;
#1 $display("%b", po);
# 1  pi=24'b110010010100001111101110;
#1 $display("%b", po);
# 1  pi=24'b101011001100010101000111;
#1 $display("%b", po);
# 1  pi=24'b001010111100111111100101;
#1 $display("%b", po);
# 1  pi=24'b000000100011010001111110;
#1 $display("%b", po);
# 1  pi=24'b010000001101011000110001;
#1 $display("%b", po);
# 1  pi=24'b100101010101111011001010;
#1 $display("%b", po);
# 1  pi=24'b011000000001011000011101;
#1 $display("%b", po);
# 1  pi=24'b001100100111111100110111;
#1 $display("%b", po);
# 1  pi=24'b100010100010010100000110;
#1 $display("%b", po);
# 1  pi=24'b111010101000100100011010;
#1 $display("%b", po);
# 1  pi=24'b001000110111111101111011;
#1 $display("%b", po);
# 1  pi=24'b100110110001001001010010;
#1 $display("%b", po);
# 1  pi=24'b001111011101111011100001;
#1 $display("%b", po);
# 1  pi=24'b101000000010010111110010;
#1 $display("%b", po);
# 1  pi=24'b011110101111011100001111;
#1 $display("%b", po);
# 1  pi=24'b110011100110000010011111;
#1 $display("%b", po);
# 1  pi=24'b101010110111010111011001;
#1 $display("%b", po);
# 1  pi=24'b100101100111111011001100;
#1 $display("%b", po);
# 1  pi=24'b001110001000011100110111;
#1 $display("%b", po);
# 1  pi=24'b111110010001010111000101;
#1 $display("%b", po);
# 1  pi=24'b011011011010011001001000;
#1 $display("%b", po);
# 1  pi=24'b000110100010000011100111;
#1 $display("%b", po);
# 1  pi=24'b110011011011011111110001;
#1 $display("%b", po);
# 1  pi=24'b011010000001100110000111;
#1 $display("%b", po);
# 1  pi=24'b000101001011110111011001;
#1 $display("%b", po);
# 1  pi=24'b110001101010110000010110;
#1 $display("%b", po);
# 1  pi=24'b110001001101101011110001;
#1 $display("%b", po);
# 1  pi=24'b110100001110010101110001;
#1 $display("%b", po);
# 1  pi=24'b001011001101011001010001;
#1 $display("%b", po);
# 1  pi=24'b000110000100011110101010;
#1 $display("%b", po);
# 1  pi=24'b011000110010110111001001;
#1 $display("%b", po);
# 1  pi=24'b100110101111110011001110;
#1 $display("%b", po);
# 1  pi=24'b000001101111101101000010;
#1 $display("%b", po);
# 1  pi=24'b001011101000100101100011;
#1 $display("%b", po);
# 1  pi=24'b111010011110111111001111;
#1 $display("%b", po);
# 1  pi=24'b001011010011100111101001;
#1 $display("%b", po);
# 1  pi=24'b111001001100110111111100;
#1 $display("%b", po);
# 1  pi=24'b001100100010000101100100;
#1 $display("%b", po);
# 1  pi=24'b010100001110100110100110;
#1 $display("%b", po);
# 1  pi=24'b011010010001000001010100;
#1 $display("%b", po);
# 1  pi=24'b001011011101110101111111;
#1 $display("%b", po);
# 1  pi=24'b001111101001011001100111;
#1 $display("%b", po);
# 1  pi=24'b001101010010011010111011;
#1 $display("%b", po);
# 1  pi=24'b001111010010111010101101;
#1 $display("%b", po);
# 1  pi=24'b010111001001100011101111;
#1 $display("%b", po);
# 1  pi=24'b011011001100010101010100;
#1 $display("%b", po);
# 1  pi=24'b000000000000100100111011;
#1 $display("%b", po);
# 1  pi=24'b100111110011101110010100;
#1 $display("%b", po);
# 1  pi=24'b011101011000111001001100;
#1 $display("%b", po);
# 1  pi=24'b010100100101100010011100;
#1 $display("%b", po);
# 1  pi=24'b101000111101001011001011;
#1 $display("%b", po);
# 1  pi=24'b010111001101100010001010;
#1 $display("%b", po);
# 1  pi=24'b100001111110101011111000;
#1 $display("%b", po);
# 1  pi=24'b000100101111010001100111;
#1 $display("%b", po);
# 1  pi=24'b111000001000001000010111;
#1 $display("%b", po);
# 1  pi=24'b011101110101000000111111;
#1 $display("%b", po);
# 1  pi=24'b100000000000111001100101;
#1 $display("%b", po);
# 1  pi=24'b001100111001001011110111;
#1 $display("%b", po);
# 1  pi=24'b110011100100010110100001;
#1 $display("%b", po);
# 1  pi=24'b001110111010101011100000;
#1 $display("%b", po);
# 1  pi=24'b000001010111010111001111;
#1 $display("%b", po);
# 1  pi=24'b000100001100000101010011;
#1 $display("%b", po);
# 1  pi=24'b000111000110101000011000;
#1 $display("%b", po);
# 1  pi=24'b101010011000000001100101;
#1 $display("%b", po);
# 1  pi=24'b100100011101000100110110;
#1 $display("%b", po);
# 1  pi=24'b001001110100011010100001;
#1 $display("%b", po);
# 1  pi=24'b101011111010100100111001;
#1 $display("%b", po);
# 1  pi=24'b010001010100000001000011;
#1 $display("%b", po);
# 1  pi=24'b011000100000111110001010;
#1 $display("%b", po);
# 1  pi=24'b000011000010111010011000;
#1 $display("%b", po);
# 1  pi=24'b011000011100101110001101;
#1 $display("%b", po);
# 1  pi=24'b100010100110101010000001;
#1 $display("%b", po);
# 1  pi=24'b010010000110100111100101;
#1 $display("%b", po);
# 1  pi=24'b110001001010001101101101;
#1 $display("%b", po);
# 1  pi=24'b001110100010101111010100;
#1 $display("%b", po);
# 1  pi=24'b001100101011111010100001;
#1 $display("%b", po);
# 1  pi=24'b100011110110100111100011;
#1 $display("%b", po);
# 1  pi=24'b011000001001111010010001;
#1 $display("%b", po);
# 1  pi=24'b110000111100000110010001;
#1 $display("%b", po);
# 1  pi=24'b001110110111110101001001;
#1 $display("%b", po);
# 1  pi=24'b011110111010111001110000;
#1 $display("%b", po);
# 1  pi=24'b010111001111010110000110;
#1 $display("%b", po);
# 1  pi=24'b000110010100011111001000;
#1 $display("%b", po);
# 1  pi=24'b011110111011101000000110;
#1 $display("%b", po);
# 1  pi=24'b111011001010101110101101;
#1 $display("%b", po);
# 1  pi=24'b010011101010101111011011;
#1 $display("%b", po);
# 1  pi=24'b111111010011101011101010;
#1 $display("%b", po);
# 1  pi=24'b100011101000011101011000;
#1 $display("%b", po);
# 1  pi=24'b001000001100001111101111;
#1 $display("%b", po);
# 1  pi=24'b000001011101100011110110;
#1 $display("%b", po);
# 1  pi=24'b100010111011000110100000;
#1 $display("%b", po);
# 1  pi=24'b111110101110111101110101;
#1 $display("%b", po);
# 1  pi=24'b000010010101100010011100;
#1 $display("%b", po);
# 1  pi=24'b011111100000010100100011;
#1 $display("%b", po);
# 1  pi=24'b110101111010010110100001;
#1 $display("%b", po);
# 1  pi=24'b100001011101011010101010;
#1 $display("%b", po);
# 1  pi=24'b000101010000011001111001;
#1 $display("%b", po);
# 1  pi=24'b101110110110000001010000;
#1 $display("%b", po);
# 1  pi=24'b100010101001100100000001;
#1 $display("%b", po);
# 1  pi=24'b001110001101110111110101;
#1 $display("%b", po);
# 1  pi=24'b100010110001011011101001;
#1 $display("%b", po);
# 1  pi=24'b001100000011001100000100;
#1 $display("%b", po);
# 1  pi=24'b111001111011101001110100;
#1 $display("%b", po);
# 1  pi=24'b001011010110111100011011;
#1 $display("%b", po);
# 1  pi=24'b011110001110101110111010;
#1 $display("%b", po);
# 1  pi=24'b100101001000110011101110;
#1 $display("%b", po);
# 1  pi=24'b011111010110010001111111;
#1 $display("%b", po);
# 1  pi=24'b010000110111011000111010;
#1 $display("%b", po);
# 1  pi=24'b100111000101011000000101;
#1 $display("%b", po);
# 1  pi=24'b001011011011111011110010;
#1 $display("%b", po);
# 1  pi=24'b111111011010000010111001;
#1 $display("%b", po);
# 1  pi=24'b000110100000110110011010;
#1 $display("%b", po);
# 1  pi=24'b011100100110101010100011;
#1 $display("%b", po);
# 1  pi=24'b111011110001100000101111;
#1 $display("%b", po);
# 1  pi=24'b110000100010110101010110;
#1 $display("%b", po);
# 1  pi=24'b110010111101101010101100;
#1 $display("%b", po);
# 1  pi=24'b111010010011000101100001;
#1 $display("%b", po);
# 1  pi=24'b100110111010001101000010;
#1 $display("%b", po);
# 1  pi=24'b101001001010010000110100;
#1 $display("%b", po);
# 1  pi=24'b011110100000100100111001;
#1 $display("%b", po);
# 1  pi=24'b001011111110011001001111;
#1 $display("%b", po);
# 1  pi=24'b111101111110111110101100;
#1 $display("%b", po);
# 1  pi=24'b011101110111011001011011;
#1 $display("%b", po);
# 1  pi=24'b001111011111010100001101;
#1 $display("%b", po);
# 1  pi=24'b011010000110101001001111;
#1 $display("%b", po);
# 1  pi=24'b111101010111100000101101;
#1 $display("%b", po);
# 1  pi=24'b101101100100011111111101;
#1 $display("%b", po);
# 1  pi=24'b111111011010110010110010;
#1 $display("%b", po);
# 1  pi=24'b010010110101001111001011;
#1 $display("%b", po);
# 1  pi=24'b010000110111101111111011;
#1 $display("%b", po);
# 1  pi=24'b111100000001000000111000;
#1 $display("%b", po);
# 1  pi=24'b000000111100100000100101;
#1 $display("%b", po);
# 1  pi=24'b000010001011110000101001;
#1 $display("%b", po);
# 1  pi=24'b010010001110101011011001;
#1 $display("%b", po);
# 1  pi=24'b101110011001100101101101;
#1 $display("%b", po);
# 1  pi=24'b101011110010100110111100;
#1 $display("%b", po);
# 1  pi=24'b010011100101101010111100;
#1 $display("%b", po);
# 1  pi=24'b011101111011000001010101;
#1 $display("%b", po);
# 1  pi=24'b111011110101011101100101;
#1 $display("%b", po);
# 1  pi=24'b001101101000111100110001;
#1 $display("%b", po);
# 1  pi=24'b101100001011101111111101;
#1 $display("%b", po);
# 1  pi=24'b001100110011011011001111;
#1 $display("%b", po);
# 1  pi=24'b001100011100000000010011;
#1 $display("%b", po);
# 1  pi=24'b010110111010111000110110;
#1 $display("%b", po);
# 1  pi=24'b100010111011011100100101;
#1 $display("%b", po);
# 1  pi=24'b001101111011001111010111;
#1 $display("%b", po);
# 1  pi=24'b011101100011100011000101;
#1 $display("%b", po);
# 1  pi=24'b010100010001111010000000;
#1 $display("%b", po);
# 1  pi=24'b010111100000000000101001;
#1 $display("%b", po);
# 1  pi=24'b101011001111100100000111;
#1 $display("%b", po);
# 1  pi=24'b100001000001100101111010;
#1 $display("%b", po);
# 1  pi=24'b100011100010010101110011;
#1 $display("%b", po);
# 1  pi=24'b110000000101110001110101;
#1 $display("%b", po);
# 1  pi=24'b110000000010110110010011;
#1 $display("%b", po);
# 1  pi=24'b011001011101110100011010;
#1 $display("%b", po);
# 1  pi=24'b011001000110011000001101;
#1 $display("%b", po);
# 1  pi=24'b001011111100001010110001;
#1 $display("%b", po);
# 1  pi=24'b010110011011010000001110;
#1 $display("%b", po);
# 1  pi=24'b001100001100100000011000;
#1 $display("%b", po);
# 1  pi=24'b000001000101010101001010;
#1 $display("%b", po);
# 1  pi=24'b101100101110110011011100;
#1 $display("%b", po);
# 1  pi=24'b100010011110011111000101;
#1 $display("%b", po);
# 1  pi=24'b101111111001011001111000;
#1 $display("%b", po);
# 1  pi=24'b110000100001010000111111;
#1 $display("%b", po);
# 1  pi=24'b000101001101100010011010;
#1 $display("%b", po);
# 1  pi=24'b011100101111101110010011;
#1 $display("%b", po);
# 1  pi=24'b111000001101111100011100;
#1 $display("%b", po);
# 1  pi=24'b000010101101011111011001;
#1 $display("%b", po);
# 1  pi=24'b111100010011100011110111;
#1 $display("%b", po);
# 1  pi=24'b101000001101011100111110;
#1 $display("%b", po);
# 1  pi=24'b001000111100101000111111;
#1 $display("%b", po);
# 1  pi=24'b010110011100000010101010;
#1 $display("%b", po);
# 1  pi=24'b110111101101101001111001;
#1 $display("%b", po);
# 1  pi=24'b011011101111110110011111;
#1 $display("%b", po);
# 1  pi=24'b011011001011111110011101;
#1 $display("%b", po);
# 1  pi=24'b101111000000001101110110;
#1 $display("%b", po);
# 1  pi=24'b101010000100100101000011;
#1 $display("%b", po);
# 1  pi=24'b100110011011000110010100;
#1 $display("%b", po);
# 1  pi=24'b000110101001011101001111;
#1 $display("%b", po);
# 1  pi=24'b100010111100011010110010;
#1 $display("%b", po);
# 1  pi=24'b110100110010000100100110;
#1 $display("%b", po);
# 1  pi=24'b111011011101011000110101;
#1 $display("%b", po);
# 1  pi=24'b001101011110010111001000;
#1 $display("%b", po);
# 1  pi=24'b010000101100010110110010;
#1 $display("%b", po);
# 1  pi=24'b010011100111011010000110;
#1 $display("%b", po);
# 1  pi=24'b101001110100111000101000;
#1 $display("%b", po);
# 1  pi=24'b001101011101000010010011;
#1 $display("%b", po);
# 1  pi=24'b111000000000011100100100;
#1 $display("%b", po);
# 1  pi=24'b101100111101101110110111;
#1 $display("%b", po);
# 1  pi=24'b100000101110110010001101;
#1 $display("%b", po);
# 1  pi=24'b110000011010111011010000;
#1 $display("%b", po);
# 1  pi=24'b001100001011100111001010;
#1 $display("%b", po);
# 1  pi=24'b110001110010110011010101;
#1 $display("%b", po);
# 1  pi=24'b010101100100101010111100;
#1 $display("%b", po);
# 1  pi=24'b000101110000110111101110;
#1 $display("%b", po);
# 1  pi=24'b001001000010110000011111;
#1 $display("%b", po);
# 1  pi=24'b010010000100100111000000;
#1 $display("%b", po);
# 1  pi=24'b000110000001110010010100;
#1 $display("%b", po);
# 1  pi=24'b011010111101100111111100;
#1 $display("%b", po);
# 1  pi=24'b011011001010110111001100;
#1 $display("%b", po);
# 1  pi=24'b101101111010111011000010;
#1 $display("%b", po);
# 1  pi=24'b001001000001000000000101;
#1 $display("%b", po);
# 1  pi=24'b101000111110001101000111;
#1 $display("%b", po);
# 1  pi=24'b010010011001011000001011;
#1 $display("%b", po);
# 1  pi=24'b010001000100010100101111;
#1 $display("%b", po);
# 1  pi=24'b000100011001100001011010;
#1 $display("%b", po);
# 1  pi=24'b000010000110001110101001;
#1 $display("%b", po);
# 1  pi=24'b000110100111110101110111;
#1 $display("%b", po);
# 1  pi=24'b010011111111111101111111;
#1 $display("%b", po);
# 1  pi=24'b010011110000111101001000;
#1 $display("%b", po);
# 1  pi=24'b011101011010111110101111;
#1 $display("%b", po);
# 1  pi=24'b000010110000000011000000;
#1 $display("%b", po);
# 1  pi=24'b011011111011010100011011;
#1 $display("%b", po);
# 1  pi=24'b010011110011001111010100;
#1 $display("%b", po);
# 1  pi=24'b111101110110001111111001;
#1 $display("%b", po);
# 1  pi=24'b000110111010101101001110;
#1 $display("%b", po);
# 1  pi=24'b100010101010000110111101;
#1 $display("%b", po);
# 1  pi=24'b101110110110101011011110;
#1 $display("%b", po);
# 1  pi=24'b001110100001111100011001;
#1 $display("%b", po);
# 1  pi=24'b101110111000101101001100;
#1 $display("%b", po);
# 1  pi=24'b011001100101000011010111;
#1 $display("%b", po);
# 1  pi=24'b001001011001111001100110;
#1 $display("%b", po);
# 1  pi=24'b111111000100001111001000;
#1 $display("%b", po);
# 1  pi=24'b110010011110011010101101;
#1 $display("%b", po);
# 1  pi=24'b111110000100000010100001;
#1 $display("%b", po);
# 1  pi=24'b000111111101010011111111;
#1 $display("%b", po);
# 1  pi=24'b100110100101000111001101;
#1 $display("%b", po);
# 1  pi=24'b101001111110111111000000;
#1 $display("%b", po);
# 1  pi=24'b100110100101011001110110;
#1 $display("%b", po);
# 1  pi=24'b011101010000111110000001;
#1 $display("%b", po);
# 1  pi=24'b011100000011000011010011;
#1 $display("%b", po);
# 1  pi=24'b010011100111100110000101;
#1 $display("%b", po);
# 1  pi=24'b010000110000101000011011;
#1 $display("%b", po);
# 1  pi=24'b101010101101010100110011;
#1 $display("%b", po);
# 1  pi=24'b110100100000101110101111;
#1 $display("%b", po);
# 1  pi=24'b011000110110110000110110;
#1 $display("%b", po);
# 1  pi=24'b101101100100011011001100;
#1 $display("%b", po);
# 1  pi=24'b001000100111101000101111;
#1 $display("%b", po);
# 1  pi=24'b110000010110000000000001;
#1 $display("%b", po);
# 1  pi=24'b001001110101100110101110;
#1 $display("%b", po);
# 1  pi=24'b110100010100110000101100;
#1 $display("%b", po);
# 1  pi=24'b001101001110000110010001;
#1 $display("%b", po);
# 1  pi=24'b110110100110110101011000;
#1 $display("%b", po);
# 1  pi=24'b111101001000011111101011;
#1 $display("%b", po);
# 1  pi=24'b010000011011010000001100;
#1 $display("%b", po);
# 1  pi=24'b010011001100101110001111;
#1 $display("%b", po);
# 1  pi=24'b101001100110000100011011;
#1 $display("%b", po);
# 1  pi=24'b111111110110110110001101;
#1 $display("%b", po);
# 1  pi=24'b100111001101101100001111;
#1 $display("%b", po);
# 1  pi=24'b001100001111011100111000;
#1 $display("%b", po);
# 1  pi=24'b001101011110110111001111;
#1 $display("%b", po);
# 1  pi=24'b110101111110001001001000;
#1 $display("%b", po);
# 1  pi=24'b000101000110010101101010;
#1 $display("%b", po);
# 1  pi=24'b011110101101110001110101;
#1 $display("%b", po);
# 1  pi=24'b011100001011100101100011;
#1 $display("%b", po);
# 1  pi=24'b010000101100100011000110;
#1 $display("%b", po);
# 1  pi=24'b001010011011000010110010;
#1 $display("%b", po);
# 1  pi=24'b000101001001011011010000;
#1 $display("%b", po);
# 1  pi=24'b000010010011011011100011;
#1 $display("%b", po);
# 1  pi=24'b011011011000110101011010;
#1 $display("%b", po);
# 1  pi=24'b001110001010101110111001;
#1 $display("%b", po);
# 1  pi=24'b011101101110111000111001;
#1 $display("%b", po);
# 1  pi=24'b111010000100000100111101;
#1 $display("%b", po);
# 1  pi=24'b001101010101000011000011;
#1 $display("%b", po);
# 1  pi=24'b001111111101001011010100;
#1 $display("%b", po);
# 1  pi=24'b111011010000000100010101;
#1 $display("%b", po);
# 1  pi=24'b100110011111101110111000;
#1 $display("%b", po);
# 1  pi=24'b100010101101011011100001;
#1 $display("%b", po);
# 1  pi=24'b101111100101111110101111;
#1 $display("%b", po);
# 1  pi=24'b111010100110110011101010;
#1 $display("%b", po);
# 1  pi=24'b011000111101011111111101;
#1 $display("%b", po);
# 1  pi=24'b001001010001000101101000;
#1 $display("%b", po);
# 1  pi=24'b000101001000000101001110;
#1 $display("%b", po);
# 1  pi=24'b001100011011110001111110;
#1 $display("%b", po);
# 1  pi=24'b001110100010100010101101;
#1 $display("%b", po);
# 1  pi=24'b001011111001100100000110;
#1 $display("%b", po);
# 1  pi=24'b011110001111111001000111;
#1 $display("%b", po);
# 1  pi=24'b110011110111010100010000;
#1 $display("%b", po);
# 1  pi=24'b001111000110101010010001;
#1 $display("%b", po);
# 1  pi=24'b000000000100100111011101;
#1 $display("%b", po);
# 1  pi=24'b011010001001111010010100;
#1 $display("%b", po);
# 1  pi=24'b110010011000100110110011;
#1 $display("%b", po);
# 1  pi=24'b110111110010101110110011;
#1 $display("%b", po);
# 1  pi=24'b000010101110000110000000;
#1 $display("%b", po);
# 1  pi=24'b000001101001000000010111;
#1 $display("%b", po);
# 1  pi=24'b101000111011110000000100;
#1 $display("%b", po);
# 1  pi=24'b111000111010111110111011;
#1 $display("%b", po);
# 1  pi=24'b001111100010010010000001;
#1 $display("%b", po);
# 1  pi=24'b111001010110010101100110;
#1 $display("%b", po);
# 1  pi=24'b110100011001111100100111;
#1 $display("%b", po);
# 1  pi=24'b011100011111111000011001;
#1 $display("%b", po);
# 1  pi=24'b011100010110110101010111;
#1 $display("%b", po);
# 1  pi=24'b000000011001111001011110;
#1 $display("%b", po);
# 1  pi=24'b110110001000000101111100;
#1 $display("%b", po);
# 1  pi=24'b111001010010100011110010;
#1 $display("%b", po);
# 1  pi=24'b111110000000111011001011;
#1 $display("%b", po);
# 1  pi=24'b100110010010101110101000;
#1 $display("%b", po);
# 1  pi=24'b101011100010010100010101;
#1 $display("%b", po);
# 1  pi=24'b010100111100110010010001;
#1 $display("%b", po);
# 1  pi=24'b001011000001101110110101;
#1 $display("%b", po);
# 1  pi=24'b111010010110111000000010;
#1 $display("%b", po);
# 1  pi=24'b110100101011100111010110;
#1 $display("%b", po);
# 1  pi=24'b011111110110101101010000;
#1 $display("%b", po);
# 1  pi=24'b101110001101011100111000;
#1 $display("%b", po);
# 1  pi=24'b001111100110111001110101;
#1 $display("%b", po);
# 1  pi=24'b110110101100000001101111;
#1 $display("%b", po);
# 1  pi=24'b000010011110111101110011;
#1 $display("%b", po);
# 1  pi=24'b001101101011111110100001;
#1 $display("%b", po);
# 1  pi=24'b101110101001010111010010;
#1 $display("%b", po);
# 1  pi=24'b111001011111100111000101;
#1 $display("%b", po);
# 1  pi=24'b110000011111100011010100;
#1 $display("%b", po);
# 1  pi=24'b010000001000111000111011;
#1 $display("%b", po);
# 1  pi=24'b100101001011010010010011;
#1 $display("%b", po);
# 1  pi=24'b010100111100010101101101;
#1 $display("%b", po);
# 1  pi=24'b100110011011111010101101;
#1 $display("%b", po);
# 1  pi=24'b110010001110111011000110;
#1 $display("%b", po);
# 1  pi=24'b010111110000101010000011;
#1 $display("%b", po);
# 1  pi=24'b010100010001001011010000;
#1 $display("%b", po);
# 1  pi=24'b010101100011010000000011;
#1 $display("%b", po);
# 1  pi=24'b001100111110111111001101;
#1 $display("%b", po);
# 1  pi=24'b110101100101000101100011;
#1 $display("%b", po);
# 1  pi=24'b111000110100000011001110;
#1 $display("%b", po);
# 1  pi=24'b000011111000011000001100;
#1 $display("%b", po);
# 1  pi=24'b010110000000000011010100;
#1 $display("%b", po);
# 1  pi=24'b100110100000110101101010;
#1 $display("%b", po);
# 1  pi=24'b011100010100101101110000;
#1 $display("%b", po);
# 1  pi=24'b011011100100110111101100;
#1 $display("%b", po);
# 1  pi=24'b101010110110001100110000;
#1 $display("%b", po);
# 1  pi=24'b001011011000010010001001;
#1 $display("%b", po);
# 1  pi=24'b000001001100001001000100;
#1 $display("%b", po);
# 1  pi=24'b110001111110100100010011;
#1 $display("%b", po);
# 1  pi=24'b100110001101101110100011;
#1 $display("%b", po);
# 1  pi=24'b010000000110111110111001;
#1 $display("%b", po);
# 1  pi=24'b100000011001110000001111;
#1 $display("%b", po);
# 1  pi=24'b011110111011100111000110;
#1 $display("%b", po);
# 1  pi=24'b011000011111110101101101;
#1 $display("%b", po);
# 1  pi=24'b100010101001000100111100;
#1 $display("%b", po);
# 1  pi=24'b001111000000010000110110;
#1 $display("%b", po);
# 1  pi=24'b110101110000010011111011;
#1 $display("%b", po);
# 1  pi=24'b111001001001000011001011;
#1 $display("%b", po);
# 1  pi=24'b110100100010010111011101;
#1 $display("%b", po);
# 1  pi=24'b010111001010111011001001;
#1 $display("%b", po);
# 1  pi=24'b110001010010111100011000;
#1 $display("%b", po);
# 1  pi=24'b001100010011110011101110;
#1 $display("%b", po);
# 1  pi=24'b010011100001011010010011;
#1 $display("%b", po);
# 1  pi=24'b000101110101111010000010;
#1 $display("%b", po);
# 1  pi=24'b111010010101001011100101;
#1 $display("%b", po);
# 1  pi=24'b001100011000101001001010;
#1 $display("%b", po);
# 1  pi=24'b010100110110000110110100;
#1 $display("%b", po);
# 1  pi=24'b001101001111110111011010;
#1 $display("%b", po);
# 1  pi=24'b100110110101010100001100;
#1 $display("%b", po);
# 1  pi=24'b001101000011010100011100;
#1 $display("%b", po);
# 1  pi=24'b000101001001000011100011;
#1 $display("%b", po);
# 1  pi=24'b010101000110111001111111;
#1 $display("%b", po);
# 1  pi=24'b000011011110011111111101;
#1 $display("%b", po);
# 1  pi=24'b011110000110011110101010;
#1 $display("%b", po);
# 1  pi=24'b001111110101001001011010;
#1 $display("%b", po);
# 1  pi=24'b010011110111011011010011;
#1 $display("%b", po);
# 1  pi=24'b100010000011100100101100;
#1 $display("%b", po);
# 1  pi=24'b101011111110111011110000;
#1 $display("%b", po);
# 1  pi=24'b110111010010100110000010;
#1 $display("%b", po);
# 1  pi=24'b101111111001110111111111;
#1 $display("%b", po);
# 1  pi=24'b010101111010000001101010;
#1 $display("%b", po);
# 1  pi=24'b001111000110001110110110;
#1 $display("%b", po);
# 1  pi=24'b010111110010101000100110;
#1 $display("%b", po);
# 1  pi=24'b100100101010001100010110;
#1 $display("%b", po);
# 1  pi=24'b001111000110111100000100;
#1 $display("%b", po);
# 1  pi=24'b101000011101011001010000;
#1 $display("%b", po);
# 1  pi=24'b111101011000010100101100;
#1 $display("%b", po);
# 1  pi=24'b011011010101110110100001;
#1 $display("%b", po);
# 1  pi=24'b010101110111101101011000;
#1 $display("%b", po);
# 1  pi=24'b010010100110001111001011;
#1 $display("%b", po);
# 1  pi=24'b111001100010010011000011;
#1 $display("%b", po);
# 1  pi=24'b101001001111000100111010;
#1 $display("%b", po);
# 1  pi=24'b001111010100011011101000;
#1 $display("%b", po);
# 1  pi=24'b001110100111101000000010;
#1 $display("%b", po);
# 1  pi=24'b010011010000110000011101;
#1 $display("%b", po);
# 1  pi=24'b100001111000100001110000;
#1 $display("%b", po);
# 1  pi=24'b100010101111110110101000;
#1 $display("%b", po);
# 1  pi=24'b110010010000000000010000;
#1 $display("%b", po);
# 1  pi=24'b000100010101010101101100;
#1 $display("%b", po);
# 1  pi=24'b000010100101010010001101;
#1 $display("%b", po);
# 1  pi=24'b010000110001100111001000;
#1 $display("%b", po);
# 1  pi=24'b010101101010011110110001;
#1 $display("%b", po);
# 1  pi=24'b111011000010100010111001;
#1 $display("%b", po);
# 1  pi=24'b001011101011100100000001;
#1 $display("%b", po);
# 1  pi=24'b101101111001101000000010;
#1 $display("%b", po);
# 1  pi=24'b011011001111000101111110;
#1 $display("%b", po);
# 1  pi=24'b100010001010100101000010;
#1 $display("%b", po);
# 1  pi=24'b001101011001010110111110;
#1 $display("%b", po);
# 1  pi=24'b011011010010101001010011;
#1 $display("%b", po);
# 1  pi=24'b110011000111110110111010;
#1 $display("%b", po);
# 1  pi=24'b101100010001110000100011;
#1 $display("%b", po);
# 1  pi=24'b110100111001001010010101;
#1 $display("%b", po);
# 1  pi=24'b000010111010001110101101;
#1 $display("%b", po);
# 1  pi=24'b100110001011001100100110;
#1 $display("%b", po);
# 1  pi=24'b010001001001110101011101;
#1 $display("%b", po);
# 1  pi=24'b110100111111000010111100;
#1 $display("%b", po);
# 1  pi=24'b100101011010000000001101;
#1 $display("%b", po);
# 1  pi=24'b011101101010011110010110;
#1 $display("%b", po);
# 1  pi=24'b010011001111001010111110;
#1 $display("%b", po);
# 1  pi=24'b010010111110000011101010;
#1 $display("%b", po);
# 1  pi=24'b110000101010000011000000;
#1 $display("%b", po);
# 1  pi=24'b001010000100110100010111;
#1 $display("%b", po);
# 1  pi=24'b101011100111100010110011;
#1 $display("%b", po);
# 1  pi=24'b001000001011101101100001;
#1 $display("%b", po);
# 1  pi=24'b111010011110010001010110;
#1 $display("%b", po);
# 1  pi=24'b010010110110000101010100;
#1 $display("%b", po);
# 1  pi=24'b011110101000111001110110;
#1 $display("%b", po);
# 1  pi=24'b110110001010010010001111;
#1 $display("%b", po);
# 1  pi=24'b111110011010111011111001;
#1 $display("%b", po);
# 1  pi=24'b101010000100011001010100;
#1 $display("%b", po);
# 1  pi=24'b110000011110001011100010;
#1 $display("%b", po);
# 1  pi=24'b011110111100011111100110;
#1 $display("%b", po);
# 1  pi=24'b110001100010010001010100;
#1 $display("%b", po);
# 1  pi=24'b100111110000010110001100;
#1 $display("%b", po);
# 1  pi=24'b100000110001000100110011;
#1 $display("%b", po);
# 1  pi=24'b001011011011011111100110;
#1 $display("%b", po);
# 1  pi=24'b110000101001100011111011;
#1 $display("%b", po);
# 1  pi=24'b100011111101110100100110;
#1 $display("%b", po);
# 1  pi=24'b111010001010100111110111;
#1 $display("%b", po);
# 1  pi=24'b100100011001101110110111;
#1 $display("%b", po);
# 1  pi=24'b010001111111011010010110;
#1 $display("%b", po);
# 1  pi=24'b111110001011000011110100;
#1 $display("%b", po);
# 1  pi=24'b100011111111011011010110;
#1 $display("%b", po);
# 1  pi=24'b001110111110111110010000;
#1 $display("%b", po);
# 1  pi=24'b110110000110000101100110;
#1 $display("%b", po);
# 1  pi=24'b011000111000011110011111;
#1 $display("%b", po);
# 1  pi=24'b100010100010011000011100;
#1 $display("%b", po);
# 1  pi=24'b011011111001000001101000;
#1 $display("%b", po);
# 1  pi=24'b100011101011100001011000;
#1 $display("%b", po);
# 1  pi=24'b101010111010110011101001;
#1 $display("%b", po);
# 1  pi=24'b101111110011010010110001;
#1 $display("%b", po);
# 1  pi=24'b011000110101101000011001;
#1 $display("%b", po);
# 1  pi=24'b001101000101110101011001;
#1 $display("%b", po);
# 1  pi=24'b101000001001111111010011;
#1 $display("%b", po);
# 1  pi=24'b111100100000111001101101;
#1 $display("%b", po);
# 1  pi=24'b100110111111111100001001;
#1 $display("%b", po);
# 1  pi=24'b001111100101101111101010;
#1 $display("%b", po);
# 1  pi=24'b111111010100011101010001;
#1 $display("%b", po);
# 1  pi=24'b010011100110011001111010;
#1 $display("%b", po);
# 1  pi=24'b111000010001010011111111;
#1 $display("%b", po);
# 1  pi=24'b100011110010101010100110;
#1 $display("%b", po);
# 1  pi=24'b000111111001101001101111;
#1 $display("%b", po);
# 1  pi=24'b000000010001011101101010;
#1 $display("%b", po);
# 1  pi=24'b101101001010110000101001;
#1 $display("%b", po);
# 1  pi=24'b110001110000100111011100;
#1 $display("%b", po);
# 1  pi=24'b011100101101101011001100;
#1 $display("%b", po);
# 1  pi=24'b000011110111111101011101;
#1 $display("%b", po);
# 1  pi=24'b001001110011111000111001;
#1 $display("%b", po);
# 1  pi=24'b001111010010111110010010;
#1 $display("%b", po);
# 1  pi=24'b011010101100110001100100;
#1 $display("%b", po);
# 1  pi=24'b000011000110011101011011;
#1 $display("%b", po);
# 1  pi=24'b110101111111011101111110;
#1 $display("%b", po);
# 1  pi=24'b110001101000111011000001;
#1 $display("%b", po);
# 1  pi=24'b000100011000011001000010;
#1 $display("%b", po);
# 1  pi=24'b011000111111100011100110;
#1 $display("%b", po);
# 1  pi=24'b110110101100101001001110;
#1 $display("%b", po);
# 1  pi=24'b100011111101100111110001;
#1 $display("%b", po);
# 1  pi=24'b000010101101101000110110;
#1 $display("%b", po);
# 1  pi=24'b111111101000010001111001;
#1 $display("%b", po);
# 1  pi=24'b011110100011010000101011;
#1 $display("%b", po);
# 1  pi=24'b100000010011110101101000;
#1 $display("%b", po);
# 1  pi=24'b010100110001100000101100;
#1 $display("%b", po);
# 1  pi=24'b100100101011101110001001;
#1 $display("%b", po);
# 1  pi=24'b101101111110011110001111;
#1 $display("%b", po);
# 1  pi=24'b100010010101111111001111;
#1 $display("%b", po);
# 1  pi=24'b101001100001010010001010;
#1 $display("%b", po);
# 1  pi=24'b110001111010101011100111;
#1 $display("%b", po);
# 1  pi=24'b001100111011111100110100;
#1 $display("%b", po);
# 1  pi=24'b111111001000100101111100;
#1 $display("%b", po);
# 1  pi=24'b011111110011101011010001;
#1 $display("%b", po);
# 1  pi=24'b011000100000011111011110;
#1 $display("%b", po);
# 1  pi=24'b011011100110101101100001;
#1 $display("%b", po);
# 1  pi=24'b000010001001011101101010;
#1 $display("%b", po);
# 1  pi=24'b010000001000111100101000;
#1 $display("%b", po);
# 1  pi=24'b110010101011101010010101;
#1 $display("%b", po);
# 1  pi=24'b111101110000000000100111;
#1 $display("%b", po);
# 1  pi=24'b011110110001010010110111;
#1 $display("%b", po);
# 1  pi=24'b111101000000101000101101;
#1 $display("%b", po);
# 1  pi=24'b011000010101000001101011;
#1 $display("%b", po);
# 1  pi=24'b110001000000101011001110;
#1 $display("%b", po);
# 1  pi=24'b010011100011101110101100;
#1 $display("%b", po);
# 1  pi=24'b010110110000010111111110;
#1 $display("%b", po);
# 1  pi=24'b010100111100000110111110;
#1 $display("%b", po);
# 1  pi=24'b000011101111000000111010;
#1 $display("%b", po);
# 1  pi=24'b110001010000001111101111;
#1 $display("%b", po);
# 1  pi=24'b011010100011011110000111;
#1 $display("%b", po);
# 1  pi=24'b011100000110100101001100;
#1 $display("%b", po);
# 1  pi=24'b100011011000110101101111;
#1 $display("%b", po);
# 1  pi=24'b111000100111000100001110;
#1 $display("%b", po);
# 1  pi=24'b001111100011000101010100;
#1 $display("%b", po);
# 1  pi=24'b111011010110011011000011;
#1 $display("%b", po);
# 1  pi=24'b001001000111100011110100;
#1 $display("%b", po);
# 1  pi=24'b101111011011011110100010;
#1 $display("%b", po);
# 1  pi=24'b000111010111111010011000;
#1 $display("%b", po);
# 1  pi=24'b100100011100111111010110;
#1 $display("%b", po);
# 1  pi=24'b011000110101100011001111;
#1 $display("%b", po);
# 1  pi=24'b110110110101000110010110;
#1 $display("%b", po);
# 1  pi=24'b100111101110001010111101;
#1 $display("%b", po);
# 1  pi=24'b011101000001100010011000;
#1 $display("%b", po);
# 1  pi=24'b001011110011111100111101;
#1 $display("%b", po);
# 1  pi=24'b011100001100111100111101;
#1 $display("%b", po);
# 1  pi=24'b001111101111111101100001;
#1 $display("%b", po);
# 1  pi=24'b010100010010101011010000;
#1 $display("%b", po);
# 1  pi=24'b010001000111111101110101;
#1 $display("%b", po);
# 1  pi=24'b001000111101000101100001;
#1 $display("%b", po);
# 1  pi=24'b001011011101001011110000;
#1 $display("%b", po);
# 1  pi=24'b111011100001010010100011;
#1 $display("%b", po);
# 1  pi=24'b010010101000000111010000;
#1 $display("%b", po);
# 1  pi=24'b110010100110111111001100;
#1 $display("%b", po);
# 1  pi=24'b101000010000000110010101;
#1 $display("%b", po);
# 1  pi=24'b011100000111110001101101;
#1 $display("%b", po);
# 1  pi=24'b100100001001111111110110;
#1 $display("%b", po);
# 1  pi=24'b101011001001000011000110;
#1 $display("%b", po);
# 1  pi=24'b110111011011010000010011;
#1 $display("%b", po);
# 1  pi=24'b111010111100111111110101;
#1 $display("%b", po);
# 1  pi=24'b111010110101001010101010;
#1 $display("%b", po);
# 1  pi=24'b000010001110000110011000;
#1 $display("%b", po);
# 1  pi=24'b011010010011010001110100;
#1 $display("%b", po);
# 1  pi=24'b100101101011101010011110;
#1 $display("%b", po);
# 1  pi=24'b111001101111010101101001;
#1 $display("%b", po);
# 1  pi=24'b011111001110011100100111;
#1 $display("%b", po);
# 1  pi=24'b010100101101000001010111;
#1 $display("%b", po);
# 1  pi=24'b011101010100110011000101;
#1 $display("%b", po);
# 1  pi=24'b011000110011010010010110;
#1 $display("%b", po);
# 1  pi=24'b111101101100000100110111;
#1 $display("%b", po);
# 1  pi=24'b011110000110111000010010;
#1 $display("%b", po);
# 1  pi=24'b111001000000100101111000;
#1 $display("%b", po);
# 1  pi=24'b000010010111101100110000;
#1 $display("%b", po);
# 1  pi=24'b101110010101100110001010;
#1 $display("%b", po);
# 1  pi=24'b110110111100110010101000;
#1 $display("%b", po);
# 1  pi=24'b110101001100101110000110;
#1 $display("%b", po);
# 1  pi=24'b001010000000100001100001;
#1 $display("%b", po);
# 1  pi=24'b111010010101110011101110;
#1 $display("%b", po);
# 1  pi=24'b010101111111101000100001;
#1 $display("%b", po);
# 1  pi=24'b010011011000011101100011;
#1 $display("%b", po);
# 1  pi=24'b110000001101100111111010;
#1 $display("%b", po);
# 1  pi=24'b111011010011101011010000;
#1 $display("%b", po);
# 1  pi=24'b101110011111001010001110;
#1 $display("%b", po);
# 1  pi=24'b110101000100011011100010;
#1 $display("%b", po);
# 1  pi=24'b110110001001101101101100;
#1 $display("%b", po);
# 1  pi=24'b011111010001001100001101;
#1 $display("%b", po);
# 1  pi=24'b110000000111000101000101;
#1 $display("%b", po);
# 1  pi=24'b001100111101110010111011;
#1 $display("%b", po);
# 1  pi=24'b011111011011101101011001;
#1 $display("%b", po);
# 1  pi=24'b000111101011001101001111;
#1 $display("%b", po);
# 1  pi=24'b000101010000101000100001;
#1 $display("%b", po);
# 1  pi=24'b011110110111011101110111;
#1 $display("%b", po);
# 1  pi=24'b010010101011000111110111;
#1 $display("%b", po);
# 1  pi=24'b110110001011111010100111;
#1 $display("%b", po);
# 1  pi=24'b001101010111010110111011;
#1 $display("%b", po);
# 1  pi=24'b100101001000110111101111;
#1 $display("%b", po);
# 1  pi=24'b110101101100001011110101;
#1 $display("%b", po);
# 1  pi=24'b111000010110100001010000;
#1 $display("%b", po);
# 1  pi=24'b100001011111011010011010;
#1 $display("%b", po);
# 1  pi=24'b101111011101111101110111;
#1 $display("%b", po);
# 1  pi=24'b101101000000111110110011;
#1 $display("%b", po);
# 1  pi=24'b110110011111101000010011;
#1 $display("%b", po);
# 1  pi=24'b011111001011111100000011;
#1 $display("%b", po);
# 1  pi=24'b010101000011010101001001;
#1 $display("%b", po);
# 1  pi=24'b011000100110100000001000;
#1 $display("%b", po);
# 1  pi=24'b000111101110011011110000;
#1 $display("%b", po);
# 1  pi=24'b011101010101110000001000;
#1 $display("%b", po);
# 1  pi=24'b001001011000000011000010;
#1 $display("%b", po);
# 1  pi=24'b100001011101100010001000;
#1 $display("%b", po);
# 1  pi=24'b010110101100101000100000;
#1 $display("%b", po);
# 1  pi=24'b010000010011000000110001;
#1 $display("%b", po);
# 1  pi=24'b111001101000110101110011;
#1 $display("%b", po);
# 1  pi=24'b111001111001011001100101;
#1 $display("%b", po);
# 1  pi=24'b110110010111011011001001;
#1 $display("%b", po);
# 1  pi=24'b100010110110110000010111;
#1 $display("%b", po);
# 1  pi=24'b010011111011100001100010;
#1 $display("%b", po);
# 1  pi=24'b000000001001001111011111;
#1 $display("%b", po);
# 1  pi=24'b111100100111001111110011;
#1 $display("%b", po);
# 1  pi=24'b100111001001001101100010;
#1 $display("%b", po);
# 1  pi=24'b100001111000001111000110;
#1 $display("%b", po);
# 1  pi=24'b001111011110010111001110;
#1 $display("%b", po);
# 1  pi=24'b101110111001110001000110;
#1 $display("%b", po);
# 1  pi=24'b101110010111101010110010;
#1 $display("%b", po);
# 1  pi=24'b010111111001100110000101;
#1 $display("%b", po);
# 1  pi=24'b001110111111010010011100;
#1 $display("%b", po);
# 1  pi=24'b010100001111111001011010;
#1 $display("%b", po);
# 1  pi=24'b001100010111001000111011;
#1 $display("%b", po);
# 1  pi=24'b111101000100101000001110;
#1 $display("%b", po);
# 1  pi=24'b000101101110111011001110;
#1 $display("%b", po);
# 1  pi=24'b100110110001000100111111;
#1 $display("%b", po);
# 1  pi=24'b010010101001111101011111;
#1 $display("%b", po);
# 1  pi=24'b101001010110100101110101;
#1 $display("%b", po);
# 1  pi=24'b111010111010000110110011;
#1 $display("%b", po);
# 1  pi=24'b111001100101111010101111;
#1 $display("%b", po);
# 1  pi=24'b111100100011001010100000;
#1 $display("%b", po);
# 1  pi=24'b101010010110001101111010;
#1 $display("%b", po);
# 1  pi=24'b110100101110011101011101;
#1 $display("%b", po);
# 1  pi=24'b010110101111110111110001;
#1 $display("%b", po);
# 1  pi=24'b101110111101010011001000;
#1 $display("%b", po);
# 1  pi=24'b011011101000111011000101;
#1 $display("%b", po);
# 1  pi=24'b000010100011101000001110;
#1 $display("%b", po);
# 1  pi=24'b100011101101111110100011;
#1 $display("%b", po);
# 1  pi=24'b110111001101100100100101;
#1 $display("%b", po);
# 1  pi=24'b000001100111110010011001;
#1 $display("%b", po);
# 1  pi=24'b101010100011011011010101;
#1 $display("%b", po);
# 1  pi=24'b111111010110001011010011;
#1 $display("%b", po);
# 1  pi=24'b000111000101000101110011;
#1 $display("%b", po);
# 1  pi=24'b111110001110111100101000;
#1 $display("%b", po);
# 1  pi=24'b000010101011101011010101;
#1 $display("%b", po);
# 1  pi=24'b011111010001010101111100;
#1 $display("%b", po);
# 1  pi=24'b100110001101001111101000;
#1 $display("%b", po);
# 1  pi=24'b000101011011011110110001;
#1 $display("%b", po);
# 1  pi=24'b100000111010101010100111;
#1 $display("%b", po);
# 1  pi=24'b000111100111111000010010;
#1 $display("%b", po);
# 1  pi=24'b001111011100110000011001;
#1 $display("%b", po);
# 1  pi=24'b110001111100011011101101;
#1 $display("%b", po);
# 1  pi=24'b110100001011100011111100;
#1 $display("%b", po);
# 1  pi=24'b001101011110110001001100;
#1 $display("%b", po);
# 1  pi=24'b111111110011100100010111;
#1 $display("%b", po);
# 1  pi=24'b111111000111100000010010;
#1 $display("%b", po);
# 1  pi=24'b101100101110111000111011;
#1 $display("%b", po);
# 1  pi=24'b010110111001000000101010;
#1 $display("%b", po);
# 1  pi=24'b100101111001001110100111;
#1 $display("%b", po);
# 1  pi=24'b110111110111001111110110;
#1 $display("%b", po);
# 1  pi=24'b101001101001111010011100;
#1 $display("%b", po);
# 1  pi=24'b011011000101001100110111;
#1 $display("%b", po);
# 1  pi=24'b100011101000001000111111;
#1 $display("%b", po);
# 1  pi=24'b100010011110010011010101;
#1 $display("%b", po);
# 1  pi=24'b000001000101000110011101;
#1 $display("%b", po);
# 1  pi=24'b101101111000010001001011;
#1 $display("%b", po);
# 1  pi=24'b111010111111101001001100;
#1 $display("%b", po);
# 1  pi=24'b010111101101001011001110;
#1 $display("%b", po);
# 1  pi=24'b100100100011100111010110;
#1 $display("%b", po);
# 1  pi=24'b100101010001000011001101;
#1 $display("%b", po);
# 1  pi=24'b010111000001110000101000;
#1 $display("%b", po);
# 1  pi=24'b001010010111111111110110;
#1 $display("%b", po);
# 1  pi=24'b001010100110011000000000;
#1 $display("%b", po);
# 1  pi=24'b110001110010111111101111;
#1 $display("%b", po);
# 1  pi=24'b100000110100000111101110;
#1 $display("%b", po);
# 1  pi=24'b001101001001100001011111;
#1 $display("%b", po);
# 1  pi=24'b001100000111100000101101;
#1 $display("%b", po);
# 1  pi=24'b110010010001001010011001;
#1 $display("%b", po);
# 1  pi=24'b110011001001011111011000;
#1 $display("%b", po);
# 1  pi=24'b011100011011111101001011;
#1 $display("%b", po);
# 1  pi=24'b011011110111010101001011;
#1 $display("%b", po);
# 1  pi=24'b000000001101110011010010;
#1 $display("%b", po);
# 1  pi=24'b001010001010010011011111;
#1 $display("%b", po);
# 1  pi=24'b100111101001010010001000;
#1 $display("%b", po);
# 1  pi=24'b001101110110010011110010;
#1 $display("%b", po);
# 1  pi=24'b100110101011010001010100;
#1 $display("%b", po);
# 1  pi=24'b000001110101100010011001;
#1 $display("%b", po);
# 1  pi=24'b111010001000101110010010;
#1 $display("%b", po);
# 1  pi=24'b011110011111010010000010;
#1 $display("%b", po);
# 1  pi=24'b011011101001000101111010;
#1 $display("%b", po);
# 1  pi=24'b011011000000001101000010;
#1 $display("%b", po);
# 1  pi=24'b011010100101000101110101;
#1 $display("%b", po);
# 1  pi=24'b011110011010001111011000;
#1 $display("%b", po);
# 1  pi=24'b111101100110111011001000;
#1 $display("%b", po);
# 1  pi=24'b011110011100110111000101;
#1 $display("%b", po);
# 1  pi=24'b000010101001011001110111;
#1 $display("%b", po);
# 1  pi=24'b011011111010000101100011;
#1 $display("%b", po);
# 1  pi=24'b001001111100011011010101;
#1 $display("%b", po);
# 1  pi=24'b000010001111111010001101;
#1 $display("%b", po);
# 1  pi=24'b000011001000001010000001;
#1 $display("%b", po);
# 1  pi=24'b011101001000001110000010;
#1 $display("%b", po);
# 1  pi=24'b110010010100001110100001;
#1 $display("%b", po);
# 1  pi=24'b100010101010100111001010;
#1 $display("%b", po);
# 1  pi=24'b000101111000100101111100;
#1 $display("%b", po);
# 1  pi=24'b011111101000111011010111;
#1 $display("%b", po);
# 1  pi=24'b100011010000111101101010;
#1 $display("%b", po);
# 1  pi=24'b110000101001001101100110;
#1 $display("%b", po);
# 1  pi=24'b000001111001100100100101;
#1 $display("%b", po);
# 1  pi=24'b111100011100101100111010;
#1 $display("%b", po);
# 1  pi=24'b110100110110010001011111;
#1 $display("%b", po);
# 1  pi=24'b001111101011010110110110;
#1 $display("%b", po);
# 1  pi=24'b101000011000001111011111;
#1 $display("%b", po);
# 1  pi=24'b111010000010101000111010;
#1 $display("%b", po);
# 1  pi=24'b111111111010000100100000;
#1 $display("%b", po);
# 1  pi=24'b001100011001000010100100;
#1 $display("%b", po);
# 1  pi=24'b111110100110101111110000;
#1 $display("%b", po);
# 1  pi=24'b010010000001010110111001;
#1 $display("%b", po);
# 1  pi=24'b111111110100010011110000;
#1 $display("%b", po);
# 1  pi=24'b111010000100000111011000;
#1 $display("%b", po);
# 1  pi=24'b010010001110101100110010;
#1 $display("%b", po);
# 1  pi=24'b111010111101001100001011;
#1 $display("%b", po);
# 1  pi=24'b011101010001011101010001;
#1 $display("%b", po);
# 1  pi=24'b100101011000000100011111;
#1 $display("%b", po);
# 1  pi=24'b110110100001010000101000;
#1 $display("%b", po);
# 1  pi=24'b001010100110100011100101;
#1 $display("%b", po);
# 1  pi=24'b001000100001011111011100;
#1 $display("%b", po);
# 1  pi=24'b100000011010110000011010;
#1 $display("%b", po);
# 1  pi=24'b011001010001100011111100;
#1 $display("%b", po);
# 1  pi=24'b001100010010110101110000;
#1 $display("%b", po);
# 1  pi=24'b011110111100010010010011;
#1 $display("%b", po);
# 1  pi=24'b001001101110000000000110;
#1 $display("%b", po);
# 1  pi=24'b011010100010001101011010;
#1 $display("%b", po);
# 1  pi=24'b010010011110110100011000;
#1 $display("%b", po);
# 1  pi=24'b101010011011110100100101;
#1 $display("%b", po);
# 1  pi=24'b100101111100001010101000;
#1 $display("%b", po);
# 1  pi=24'b111100101001101010111111;
#1 $display("%b", po);
# 1  pi=24'b100110110100000011101010;
#1 $display("%b", po);
# 1  pi=24'b001100000011100011101110;
#1 $display("%b", po);
# 1  pi=24'b111011000011010101101111;
#1 $display("%b", po);
# 1  pi=24'b001100111100111010000100;
#1 $display("%b", po);
# 1  pi=24'b001000110001011010101000;
#1 $display("%b", po);
# 1  pi=24'b011111101110110101000110;
#1 $display("%b", po);
# 1  pi=24'b010011100111000010000010;
#1 $display("%b", po);
# 1  pi=24'b000011000111100011011010;
#1 $display("%b", po);
# 1  pi=24'b001100000100000000101100;
#1 $display("%b", po);
# 1  pi=24'b111110100100000010000001;
#1 $display("%b", po);
# 1  pi=24'b111001111000010110000100;
#1 $display("%b", po);
# 1  pi=24'b100000111100011111110110;
#1 $display("%b", po);
# 1  pi=24'b110000011010000000011001;
#1 $display("%b", po);
# 1  pi=24'b010100010010111011110100;
#1 $display("%b", po);
# 1  pi=24'b101010011101001000011000;
#1 $display("%b", po);
# 1  pi=24'b011000100011110001100111;
#1 $display("%b", po);
# 1  pi=24'b111010001011011011011010;
#1 $display("%b", po);
# 1  pi=24'b010111111001111000001001;
#1 $display("%b", po);
# 1  pi=24'b010010011010010001110101;
#1 $display("%b", po);
# 1  pi=24'b111111100011000001101100;
#1 $display("%b", po);
# 1  pi=24'b010001000010111100100100;
#1 $display("%b", po);
# 1  pi=24'b100010110000101100011111;
#1 $display("%b", po);
# 1  pi=24'b011100101010001001110001;
#1 $display("%b", po);
# 1  pi=24'b111101100101100011101011;
#1 $display("%b", po);
# 1  pi=24'b011011011100111010111111;
#1 $display("%b", po);
# 1  pi=24'b010100000100100000001111;
#1 $display("%b", po);
# 1  pi=24'b101101101010011110100110;
#1 $display("%b", po);
# 1  pi=24'b111011001100100110111110;
#1 $display("%b", po);
# 1  pi=24'b110011011110000100100110;
#1 $display("%b", po);
# 1  pi=24'b000010011011100001010010;
#1 $display("%b", po);
# 1  pi=24'b110000111001111011000111;
#1 $display("%b", po);
# 1  pi=24'b111011110110010011110111;
#1 $display("%b", po);
# 1  pi=24'b101011010010100100001111;
#1 $display("%b", po);
# 1  pi=24'b000000000101110110001101;
#1 $display("%b", po);
# 1  pi=24'b111001101010100111011111;
#1 $display("%b", po);
# 1  pi=24'b011100000001011111001100;
#1 $display("%b", po);
# 1  pi=24'b111110100110011110101011;
#1 $display("%b", po);
# 1  pi=24'b001000110010010101011101;
#1 $display("%b", po);
# 1  pi=24'b110100110110010000101101;
#1 $display("%b", po);
# 1  pi=24'b101000000011101011110000;
#1 $display("%b", po);
# 1  pi=24'b011101101010000111110110;
#1 $display("%b", po);
# 1  pi=24'b000110011011110101000101;
#1 $display("%b", po);
# 1  pi=24'b000000110101111110111111;
#1 $display("%b", po);
# 1  pi=24'b001001010111000101001011;
#1 $display("%b", po);
# 1  pi=24'b010100010001111101001111;
#1 $display("%b", po);
# 1  pi=24'b111111100000110110011110;
#1 $display("%b", po);
# 1  pi=24'b111011110110000100110000;
#1 $display("%b", po);
# 1  pi=24'b010000001011010010100011;
#1 $display("%b", po);
# 1  pi=24'b110101011011111111010000;
#1 $display("%b", po);
# 1  pi=24'b001011010011110101001001;
#1 $display("%b", po);
# 1  pi=24'b001000000110000111101010;
#1 $display("%b", po);
# 1  pi=24'b000111011111001100000110;
#1 $display("%b", po);
# 1  pi=24'b011001101101011000100000;
#1 $display("%b", po);
# 1  pi=24'b101001110000100110111001;
#1 $display("%b", po);
# 1  pi=24'b001001011110110101111111;
#1 $display("%b", po);
# 1  pi=24'b100011000100011101101110;
#1 $display("%b", po);
# 1  pi=24'b110111010101010100101110;
#1 $display("%b", po);
# 1  pi=24'b101100011001110001001110;
#1 $display("%b", po);
# 1  pi=24'b011100010110110111111001;
#1 $display("%b", po);
# 1  pi=24'b010110101011011110000101;
#1 $display("%b", po);
# 1  pi=24'b001110000110000100111101;
#1 $display("%b", po);
# 1  pi=24'b110000101011101010110000;
#1 $display("%b", po);
# 1  pi=24'b011111100110111100001101;
#1 $display("%b", po);
# 1  pi=24'b100100101000011101011001;
#1 $display("%b", po);
# 1  pi=24'b010000101110101101100111;
#1 $display("%b", po);
# 1  pi=24'b100110001110101011010010;
#1 $display("%b", po);
# 1  pi=24'b100101101101111100001001;
#1 $display("%b", po);
# 1  pi=24'b000111000010011101010000;
#1 $display("%b", po);
# 1  pi=24'b000100111001110010001000;
#1 $display("%b", po);
# 1  pi=24'b000000110110001100001000;
#1 $display("%b", po);
# 1  pi=24'b010000001000111010110010;
#1 $display("%b", po);
# 1  pi=24'b011000000111101111111111;
#1 $display("%b", po);
# 1  pi=24'b011101000000000010001011;
#1 $display("%b", po);
# 1  pi=24'b101110111111110100001101;
#1 $display("%b", po);
# 1  pi=24'b001011001011100011001011;
#1 $display("%b", po);
# 1  pi=24'b000100100111000000010011;
#1 $display("%b", po);
# 1  pi=24'b110000100111110011101110;
#1 $display("%b", po);
# 1  pi=24'b010011100101010010111011;
#1 $display("%b", po);
# 1  pi=24'b101000010001001111010010;
#1 $display("%b", po);
# 1  pi=24'b001001101100000000001101;
#1 $display("%b", po);
# 1  pi=24'b101000111000011000000010;
#1 $display("%b", po);
# 1  pi=24'b100011110101011010100111;
#1 $display("%b", po);
# 1  pi=24'b000101101001000001111010;
#1 $display("%b", po);
# 1  pi=24'b001000000011000001110100;
#1 $display("%b", po);
# 1  pi=24'b010010110111001011111011;
#1 $display("%b", po);
# 1  pi=24'b100000010001111001101101;
#1 $display("%b", po);
# 1  pi=24'b000010100111111011100110;
#1 $display("%b", po);
# 1  pi=24'b100010010011101000010110;
#1 $display("%b", po);
# 1  pi=24'b110110100111111110011100;
#1 $display("%b", po);
# 1  pi=24'b100010001101101001010111;
#1 $display("%b", po);
# 1  pi=24'b001001101011011110101110;
#1 $display("%b", po);
# 1  pi=24'b010010010010001011001000;
#1 $display("%b", po);
# 1  pi=24'b011100010110100010010011;
#1 $display("%b", po);
# 1  pi=24'b111101001100001111111111;
#1 $display("%b", po);
# 1  pi=24'b111111001101011001110101;
#1 $display("%b", po);
# 1  pi=24'b110010111000010010111000;
#1 $display("%b", po);
# 1  pi=24'b011110101101010001001110;
#1 $display("%b", po);
# 1  pi=24'b000101000011111000101010;
#1 $display("%b", po);
# 1  pi=24'b100000100110001111110001;
#1 $display("%b", po);
# 1  pi=24'b000010100110000110101000;
#1 $display("%b", po);
# 1  pi=24'b011101010111001101011011;
#1 $display("%b", po);
# 1  pi=24'b101010100101011011111100;
#1 $display("%b", po);
# 1  pi=24'b100111110010001110001111;
#1 $display("%b", po);
# 1  pi=24'b001011110110101110000111;
#1 $display("%b", po);
# 1  pi=24'b100101111100011110000010;
#1 $display("%b", po);
# 1  pi=24'b100011001101001010101110;
#1 $display("%b", po);
# 1  pi=24'b011001100101100000000011;
#1 $display("%b", po);
# 1  pi=24'b001010001101100111001101;
#1 $display("%b", po);
# 1  pi=24'b111100100011011010001100;
#1 $display("%b", po);
# 1  pi=24'b001110110011111111100101;
#1 $display("%b", po);
# 1  pi=24'b001010101101100101011011;
#1 $display("%b", po);
# 1  pi=24'b100100111111100100011010;
#1 $display("%b", po);
# 1  pi=24'b110010010011011010010000;
#1 $display("%b", po);
# 1  pi=24'b101100100111011010011101;
#1 $display("%b", po);
# 1  pi=24'b001110001111110101101101;
#1 $display("%b", po);
# 1  pi=24'b100110000100101111011100;
#1 $display("%b", po);
# 1  pi=24'b110001111010001110010010;
#1 $display("%b", po);
# 1  pi=24'b000000010010000001100010;
#1 $display("%b", po);
# 1  pi=24'b000111101000010110001111;
#1 $display("%b", po);
# 1  pi=24'b011111001111111001110111;
#1 $display("%b", po);
# 1  pi=24'b010110100011001000100110;
#1 $display("%b", po);
# 1  pi=24'b110011011110100001000101;
#1 $display("%b", po);
# 1  pi=24'b101101100010001001110101;
#1 $display("%b", po);
# 1  pi=24'b000001101000101011010001;
#1 $display("%b", po);
# 1  pi=24'b010011001101100010111001;
#1 $display("%b", po);
# 1  pi=24'b100110110001000111100101;
#1 $display("%b", po);
# 1  pi=24'b100001010011101110110101;
#1 $display("%b", po);
# 1  pi=24'b001010110001010110111101;
#1 $display("%b", po);
# 1  pi=24'b000000001010111001010111;
#1 $display("%b", po);
# 1  pi=24'b011110011001101100111000;
#1 $display("%b", po);
# 1  pi=24'b111111110100010000111010;
#1 $display("%b", po);
# 1  pi=24'b010000010001101111110100;
#1 $display("%b", po);
# 1  pi=24'b010001110010100110011010;
#1 $display("%b", po);
# 1  pi=24'b100011111011100000010100;
#1 $display("%b", po);
# 1  pi=24'b110001001111011101010111;
#1 $display("%b", po);
# 1  pi=24'b101000001111011110011001;
#1 $display("%b", po);
# 1  pi=24'b111111001101101011000010;
#1 $display("%b", po);
# 1  pi=24'b001001000011001111110001;
#1 $display("%b", po);
# 1  pi=24'b001110001110111010001110;
#1 $display("%b", po);
# 1  pi=24'b111000001001101111110111;
#1 $display("%b", po);
# 1  pi=24'b110001011101110100010011;
#1 $display("%b", po);
# 1  pi=24'b100000101011101011110111;
#1 $display("%b", po);
# 1  pi=24'b011000001001110110000100;
#1 $display("%b", po);
# 1  pi=24'b101010111011011001000111;
#1 $display("%b", po);
# 1  pi=24'b100110111110100100000011;
#1 $display("%b", po);
# 1  pi=24'b011100111100100001000100;
#1 $display("%b", po);
# 1  pi=24'b100000101010100111000000;
#1 $display("%b", po);
# 1  pi=24'b110001000011111100111111;
#1 $display("%b", po);
# 1  pi=24'b101100011110100101111111;
#1 $display("%b", po);
# 1  pi=24'b011011100001101011000110;
#1 $display("%b", po);
# 1  pi=24'b100100111001000101111010;
#1 $display("%b", po);
# 1  pi=24'b011001110000001110110011;
#1 $display("%b", po);
# 1  pi=24'b110101111110001001110101;
#1 $display("%b", po);
# 1  pi=24'b110001001000110000110000;
#1 $display("%b", po);
# 1  pi=24'b010101110011111010011101;
#1 $display("%b", po);
# 1  pi=24'b111001100100001001000101;
#1 $display("%b", po);
# 1  pi=24'b111110101010101111100101;
#1 $display("%b", po);
# 1  pi=24'b111001011110101111011000;
#1 $display("%b", po);
# 1  pi=24'b101000100111011100100110;
#1 $display("%b", po);
# 1  pi=24'b000001010010101000100111;
#1 $display("%b", po);
# 1  pi=24'b110111010111110011001000;
#1 $display("%b", po);
# 1  pi=24'b100101011111011011110010;
#1 $display("%b", po);
# 1  pi=24'b000100011101011101001001;
#1 $display("%b", po);
# 1  pi=24'b010110001100011101010111;
#1 $display("%b", po);
# 1  pi=24'b101100010000000110010000;
#1 $display("%b", po);
# 1  pi=24'b000111011101001110110101;
#1 $display("%b", po);
# 1  pi=24'b001010111010011101001000;
#1 $display("%b", po);
# 1  pi=24'b100001110010000101100000;
#1 $display("%b", po);
# 1  pi=24'b100100010010110100001000;
#1 $display("%b", po);
# 1  pi=24'b011101110001011100000000;
#1 $display("%b", po);
# 1  pi=24'b010011111000110110010100;
#1 $display("%b", po);
# 1  pi=24'b110111010011001001000011;
#1 $display("%b", po);
# 1  pi=24'b001111101010100111100001;
#1 $display("%b", po);
# 1  pi=24'b101010011110100010111010;
#1 $display("%b", po);
# 1  pi=24'b100110000011111011011101;
#1 $display("%b", po);
# 1  pi=24'b010101100000010000111001;
#1 $display("%b", po);
# 1  pi=24'b111101110111001100100110;
#1 $display("%b", po);
# 1  pi=24'b001011101011111110000110;
#1 $display("%b", po);
# 1  pi=24'b010010110001011110101011;
#1 $display("%b", po);
# 1  pi=24'b010010010001100000100011;
#1 $display("%b", po);
# 1  pi=24'b000100100101110110010010;
#1 $display("%b", po);
# 1  pi=24'b000110001101010100000100;
#1 $display("%b", po);
# 1  pi=24'b101011101010010001110111;
#1 $display("%b", po);
# 1  pi=24'b010001100101110111010001;
#1 $display("%b", po);
# 1  pi=24'b111110101011000111100000;
#1 $display("%b", po);
# 1  pi=24'b101110001010111100011101;
#1 $display("%b", po);
# 1  pi=24'b000101011111010100011000;
#1 $display("%b", po);
# 1  pi=24'b001011011010101111110011;
#1 $display("%b", po);
# 1  pi=24'b110010011111011001111111;
#1 $display("%b", po);
# 1  pi=24'b010011010100101111111111;
#1 $display("%b", po);
# 1  pi=24'b010100001011110001010011;
#1 $display("%b", po);
# 1  pi=24'b000101000101001010101001;
#1 $display("%b", po);
# 1  pi=24'b001100111101101000011010;
#1 $display("%b", po);
# 1  pi=24'b010000100111110101000001;
#1 $display("%b", po);
# 1  pi=24'b001010101000011110111011;
#1 $display("%b", po);
# 1  pi=24'b000110100100010000010101;
#1 $display("%b", po);
# 1  pi=24'b000000101010001011111101;
#1 $display("%b", po);
# 1  pi=24'b000000000110000011101111;
#1 $display("%b", po);
# 1  pi=24'b111001000010001011001110;
#1 $display("%b", po);
# 1  pi=24'b101100000101111100011011;
#1 $display("%b", po);
# 1  pi=24'b101110001010101010111101;
#1 $display("%b", po);
# 1  pi=24'b000101101100110110001110;
#1 $display("%b", po);
# 1  pi=24'b100011010000100110110100;
#1 $display("%b", po);
# 1  pi=24'b010110111000011000001000;
#1 $display("%b", po);
# 1  pi=24'b100101101011101010111000;
#1 $display("%b", po);
# 1  pi=24'b110000111110111111101101;
#1 $display("%b", po);
# 1  pi=24'b001100011011111110101100;
#1 $display("%b", po);
# 1  pi=24'b100011000010111110111000;
#1 $display("%b", po);
# 1  pi=24'b000001100110001011101000;
#1 $display("%b", po);
# 1  pi=24'b100110000110100000100101;
#1 $display("%b", po);
# 1  pi=24'b011101100000001111000000;
#1 $display("%b", po);
# 1  pi=24'b110001100010011101110111;
#1 $display("%b", po);
# 1  pi=24'b000000101110100101000110;
#1 $display("%b", po);
# 1  pi=24'b101101111010011100100101;
#1 $display("%b", po);
# 1  pi=24'b001100110110101100010110;
#1 $display("%b", po);
# 1  pi=24'b110010011111100100111011;
#1 $display("%b", po);
# 1  pi=24'b111001111110010011011010;
#1 $display("%b", po);
# 1  pi=24'b101100111111011110100000;
#1 $display("%b", po);
# 1  pi=24'b010010000010001010010001;
#1 $display("%b", po);
# 1  pi=24'b101011000110001110101110;
#1 $display("%b", po);
# 1  pi=24'b010010001001010000101110;
#1 $display("%b", po);
# 1  pi=24'b101101001101110000111111;
#1 $display("%b", po);
# 1  pi=24'b010010001101010010001101;
#1 $display("%b", po);
# 1  pi=24'b111000000111111011010111;
#1 $display("%b", po);
# 1  pi=24'b010011101101001001111101;
#1 $display("%b", po);
# 1  pi=24'b110011001010100111101000;
#1 $display("%b", po);
# 1  pi=24'b001001101011100110010110;
#1 $display("%b", po);
# 1  pi=24'b000001100010010001001111;
#1 $display("%b", po);
# 1  pi=24'b011001001100000011010001;
#1 $display("%b", po);
# 1  pi=24'b100100011101110100011101;
#1 $display("%b", po);
# 1  pi=24'b110100101010000011000000;
#1 $display("%b", po);
# 1  pi=24'b100111110111101100001001;
#1 $display("%b", po);
# 1  pi=24'b100011110000111010110011;
#1 $display("%b", po);
# 1  pi=24'b000011111110011000000100;
#1 $display("%b", po);
# 1  pi=24'b100100011110001001101110;
#1 $display("%b", po);
# 1  pi=24'b000101110010000001000111;
#1 $display("%b", po);
# 1  pi=24'b111010001000010000111010;
#1 $display("%b", po);
# 1  pi=24'b100001010111101101011011;
#1 $display("%b", po);
# 1  pi=24'b110101101100001101010011;
#1 $display("%b", po);
# 1  pi=24'b010111011101010001011100;
#1 $display("%b", po);
# 1  pi=24'b000010111010011110110000;
#1 $display("%b", po);
# 1  pi=24'b011110010101111111110101;
#1 $display("%b", po);
# 1  pi=24'b001100001000110001110001;
#1 $display("%b", po);
# 1  pi=24'b000001001111110110001010;
#1 $display("%b", po);
# 1  pi=24'b000101001101001110000011;
#1 $display("%b", po);
# 1  pi=24'b010100100110101110001110;
#1 $display("%b", po);
# 1  pi=24'b110101000111010100100011;
#1 $display("%b", po);
# 1  pi=24'b110011101111011010000111;
#1 $display("%b", po);
# 1  pi=24'b011100010100101111101111;
#1 $display("%b", po);
# 1  pi=24'b101111111001101000110110;
#1 $display("%b", po);
# 1  pi=24'b110110001111101011011100;
#1 $display("%b", po);
# 1  pi=24'b100011011100110101011101;
#1 $display("%b", po);
# 1  pi=24'b101110000101101000111010;
#1 $display("%b", po);
# 1  pi=24'b000010111110011111111001;
#1 $display("%b", po);
# 1  pi=24'b100000010101011110110101;
#1 $display("%b", po);
# 1  pi=24'b111011110111000110100011;
#1 $display("%b", po);
# 1  pi=24'b111001000110010111001101;
#1 $display("%b", po);
# 1  pi=24'b101011000000000110011100;
#1 $display("%b", po);
# 1  pi=24'b111011011011001010110111;
#1 $display("%b", po);
# 1  pi=24'b011000001100101011100011;
#1 $display("%b", po);
# 1  pi=24'b111111101111010100000001;
#1 $display("%b", po);
# 1  pi=24'b010010011000000011010010;
#1 $display("%b", po);
# 1  pi=24'b100001101100100100001010;
#1 $display("%b", po);
# 1  pi=24'b111000101011110010101110;
#1 $display("%b", po);
# 1  pi=24'b011011100011101010111000;
#1 $display("%b", po);
# 1  pi=24'b001010110110001111001001;
#1 $display("%b", po);
# 1  pi=24'b010101010101100100011100;
#1 $display("%b", po);
# 1  pi=24'b001010110111000101100011;
#1 $display("%b", po);
# 1  pi=24'b101111100101010101000110;
#1 $display("%b", po);
# 1  pi=24'b100000101111010110100100;
#1 $display("%b", po);
# 1  pi=24'b100101111110101110111110;
#1 $display("%b", po);
# 1  pi=24'b101100111001011010101100;
#1 $display("%b", po);
# 1  pi=24'b010111010110011010001001;
#1 $display("%b", po);
# 1  pi=24'b101000010011001110101011;
#1 $display("%b", po);
# 1  pi=24'b110001000010001011011101;
#1 $display("%b", po);
# 1  pi=24'b100111110010100101101001;
#1 $display("%b", po);
# 1  pi=24'b111011000010100100110011;
#1 $display("%b", po);
# 1  pi=24'b011010001000111011000010;
#1 $display("%b", po);
# 1  pi=24'b001101100110101011101000;
#1 $display("%b", po);
# 1  pi=24'b001011100110110101000111;
#1 $display("%b", po);
# 1  pi=24'b111011111000001010001101;
#1 $display("%b", po);
# 1  pi=24'b000100111010110100110101;
#1 $display("%b", po);
# 1  pi=24'b000010010011101010110000;
#1 $display("%b", po);
# 1  pi=24'b100000001001010100000110;
#1 $display("%b", po);
# 1  pi=24'b110110100110001011001000;
#1 $display("%b", po);
# 1  pi=24'b110100011001110011001000;
#1 $display("%b", po);
# 1  pi=24'b001111011001100000010101;
#1 $display("%b", po);
# 1  pi=24'b001000100101100011100100;
#1 $display("%b", po);
# 1  pi=24'b111011010111000011001010;
#1 $display("%b", po);
# 1  pi=24'b011101001010101101000100;
#1 $display("%b", po);
# 1  pi=24'b000110101111101010000010;
#1 $display("%b", po);
# 1  pi=24'b010100000010001010011100;
#1 $display("%b", po);
# 1  pi=24'b111000010100110111001111;
#1 $display("%b", po);
# 1  pi=24'b110101011001110010110100;
#1 $display("%b", po);
# 1  pi=24'b010101111111100000100001;
#1 $display("%b", po);
# 1  pi=24'b101011001111000001101001;
#1 $display("%b", po);
# 1  pi=24'b100001000101111011011010;
#1 $display("%b", po);
# 1  pi=24'b000101100011111111001011;
#1 $display("%b", po);
# 1  pi=24'b111111100100111101010010;
#1 $display("%b", po);
# 1  pi=24'b111001111001000100101110;
#1 $display("%b", po);
# 1  pi=24'b111011010101001110010000;
#1 $display("%b", po);
# 1  pi=24'b011000001111111011001100;
#1 $display("%b", po);
# 1  pi=24'b100110011100000110100101;
#1 $display("%b", po);
# 1  pi=24'b101001111110001000111001;
#1 $display("%b", po);
# 1  pi=24'b101000111100010110010110;
#1 $display("%b", po);
# 1  pi=24'b110111000011111101010001;
#1 $display("%b", po);
# 1  pi=24'b011000100111101011110111;
#1 $display("%b", po);
# 1  pi=24'b001100011101000100011001;
#1 $display("%b", po);
# 1  pi=24'b111111111001101110011110;
#1 $display("%b", po);
# 1  pi=24'b111110101110010101011110;
#1 $display("%b", po);
# 1  pi=24'b010000010000111111001110;
#1 $display("%b", po);
# 1  pi=24'b011001110100110001010010;
#1 $display("%b", po);
# 1  pi=24'b000101111010101000000011;
#1 $display("%b", po);
# 1  pi=24'b000010101100010011110011;
#1 $display("%b", po);
# 1  pi=24'b100000111011011101101101;
#1 $display("%b", po);
# 1  pi=24'b011001101100111010110010;
#1 $display("%b", po);
# 1  pi=24'b101001111111100000011100;
#1 $display("%b", po);
# 1  pi=24'b001000001101001010110101;
#1 $display("%b", po);
# 1  pi=24'b000011000011010010000011;
#1 $display("%b", po);
# 1  pi=24'b111110001000001110001110;
#1 $display("%b", po);
# 1  pi=24'b101101110001010010100111;
#1 $display("%b", po);
# 1  pi=24'b010100011101011000111010;
#1 $display("%b", po);
# 1  pi=24'b100011000111001110001010;
#1 $display("%b", po);
# 1  pi=24'b101010011000110101010100;
#1 $display("%b", po);
# 1  pi=24'b101000011000101111000110;
#1 $display("%b", po);
# 1  pi=24'b101011100001011110110001;
#1 $display("%b", po);
# 1  pi=24'b000111011001101100010111;
#1 $display("%b", po);
# 1  pi=24'b101001011101001001010100;
#1 $display("%b", po);
# 1  pi=24'b000010001011000011100110;
#1 $display("%b", po);
# 1  pi=24'b010000000011000101111010;
#1 $display("%b", po);
# 1  pi=24'b100010010100000110110110;
#1 $display("%b", po);
# 1  pi=24'b100010111011100100110101;
#1 $display("%b", po);
# 1  pi=24'b000100110111100010110110;
#1 $display("%b", po);
# 1  pi=24'b100010001001111101000011;
#1 $display("%b", po);
# 1  pi=24'b111000001100001100100000;
#1 $display("%b", po);
# 1  pi=24'b101111011100001001100110;
#1 $display("%b", po);
# 1  pi=24'b100101001100110000000000;
#1 $display("%b", po);
# 1  pi=24'b110010100010010011111011;
#1 $display("%b", po);
# 1  pi=24'b100100101001100001110011;
#1 $display("%b", po);
# 1  pi=24'b101000101101000110110100;
#1 $display("%b", po);
# 1  pi=24'b100111110111101110011100;
#1 $display("%b", po);
# 1  pi=24'b100000101011111111000101;
#1 $display("%b", po);
# 1  pi=24'b010100100111000010100001;
#1 $display("%b", po);
# 1  pi=24'b100110001110011110010101;
#1 $display("%b", po);
# 1  pi=24'b010100110101000000101100;
#1 $display("%b", po);
# 1  pi=24'b100100110000001001010001;
#1 $display("%b", po);
# 1  pi=24'b101010010111001101000001;
#1 $display("%b", po);
# 1  pi=24'b010100011000001010110101;
#1 $display("%b", po);
# 1  pi=24'b011000011100010001101101;
#1 $display("%b", po);
# 1  pi=24'b110100011101100100001010;
#1 $display("%b", po);
# 1  pi=24'b100010110000001000111000;
#1 $display("%b", po);
# 1  pi=24'b101010101101110101001111;
#1 $display("%b", po);
# 1  pi=24'b010100101111101101100001;
#1 $display("%b", po);
# 1  pi=24'b011101010001101110100011;
#1 $display("%b", po);
# 1  pi=24'b010101101111110001101011;
#1 $display("%b", po);
# 1  pi=24'b101000001100111010101000;
#1 $display("%b", po);
# 1  pi=24'b001101110111011011111001;
#1 $display("%b", po);
# 1  pi=24'b011101111110011010000001;
#1 $display("%b", po);
# 1  pi=24'b101101010111111101100110;
#1 $display("%b", po);
# 1  pi=24'b010110001100000101111011;
#1 $display("%b", po);
# 1  pi=24'b100000111100000010111011;
#1 $display("%b", po);
# 1  pi=24'b001100001010010110101111;
#1 $display("%b", po);
# 1  pi=24'b111101001100010000000001;
#1 $display("%b", po);
# 1  pi=24'b011010000111101001000111;
#1 $display("%b", po);
# 1  pi=24'b100101111101100111100011;
#1 $display("%b", po);
# 1  pi=24'b010011000011110001111111;
#1 $display("%b", po);
# 1  pi=24'b101011001101111000010101;
#1 $display("%b", po);
# 1  pi=24'b111101010101011100001011;
#1 $display("%b", po);
# 1  pi=24'b001100001000110111001001;
#1 $display("%b", po);
# 1  pi=24'b110000100011011100111101;
#1 $display("%b", po);
# 1  pi=24'b110001001000101100011011;
#1 $display("%b", po);
# 1  pi=24'b111110100101110101010010;
#1 $display("%b", po);
# 1  pi=24'b001001101110101000000110;
#1 $display("%b", po);
# 1  pi=24'b101111011011100110001111;
#1 $display("%b", po);
# 1  pi=24'b100000111000000111111100;
#1 $display("%b", po);
# 1  pi=24'b110111110101101101110011;
#1 $display("%b", po);
# 1  pi=24'b011111111001010111010110;
#1 $display("%b", po);
# 1  pi=24'b101000111101010111111101;
#1 $display("%b", po);
# 1  pi=24'b000111101000010101001101;
#1 $display("%b", po);
# 1  pi=24'b101110101011100111100000;
#1 $display("%b", po);
# 1  pi=24'b001110101100010111100011;
#1 $display("%b", po);
# 1  pi=24'b001111010100101000011010;
#1 $display("%b", po);
# 1  pi=24'b111011111100011110100001;
#1 $display("%b", po);
# 1  pi=24'b111000100011010111000000;
#1 $display("%b", po);
# 1  pi=24'b001101000010000011100010;
#1 $display("%b", po);
# 1  pi=24'b111110001000100000011101;
#1 $display("%b", po);
# 1  pi=24'b001110100100110011010000;
#1 $display("%b", po);
# 1  pi=24'b111101101111110100000100;
#1 $display("%b", po);
# 1  pi=24'b001001000000110110000100;
#1 $display("%b", po);
# 1  pi=24'b111011101101101101001101;
#1 $display("%b", po);
# 1  pi=24'b110100110010001011001010;
#1 $display("%b", po);
# 1  pi=24'b010000110101101111100111;
#1 $display("%b", po);
# 1  pi=24'b000011010001110110011000;
#1 $display("%b", po);
# 1  pi=24'b011001000010000111011000;
#1 $display("%b", po);
# 1  pi=24'b000101010001000000110010;
#1 $display("%b", po);
# 1  pi=24'b111110010111010001010110;
#1 $display("%b", po);
# 1  pi=24'b010100011100111111100000;
#1 $display("%b", po);
# 1  pi=24'b101110010110011001001010;
#1 $display("%b", po);
# 1  pi=24'b110001000010110100000010;
#1 $display("%b", po);
# 1  pi=24'b110100001100011100010011;
#1 $display("%b", po);
# 1  pi=24'b000011000101011010011111;
#1 $display("%b", po);
# 1  pi=24'b110111010000010111111010;
#1 $display("%b", po);
# 1  pi=24'b111100000011011011111011;
#1 $display("%b", po);
# 1  pi=24'b001010001101010111100010;
#1 $display("%b", po);
# 1  pi=24'b011111011101110100101110;
#1 $display("%b", po);
# 1  pi=24'b010110011001001101011011;
#1 $display("%b", po);
# 1  pi=24'b111000110110110000011111;
#1 $display("%b", po);
# 1  pi=24'b000101001111001101101001;
#1 $display("%b", po);
# 1  pi=24'b101110010000001100000110;
#1 $display("%b", po);
# 1  pi=24'b111111001000001111010011;
#1 $display("%b", po);
# 1  pi=24'b011010000110110110011101;
#1 $display("%b", po);
# 1  pi=24'b011101000010000001010010;
#1 $display("%b", po);
# 1  pi=24'b101101001011110111101011;
#1 $display("%b", po);
# 1  pi=24'b101111000010000000101000;
#1 $display("%b", po);
# 1  pi=24'b000010000001011001101111;
#1 $display("%b", po);
# 1  pi=24'b110101011101111000010000;
#1 $display("%b", po);
# 1  pi=24'b110001000000100111101001;
#1 $display("%b", po);
# 1  pi=24'b101111011011000001011110;
#1 $display("%b", po);
# 1  pi=24'b101100011111100010110111;
#1 $display("%b", po);
# 1  pi=24'b111111001101110000001000;
#1 $display("%b", po);
# 1  pi=24'b001001011010000001000111;
#1 $display("%b", po);
# 1  pi=24'b111110100001001010101010;
#1 $display("%b", po);
# 1  pi=24'b010001011010101010110101;
#1 $display("%b", po);
# 1  pi=24'b011001111110110001100111;
#1 $display("%b", po);
# 1  pi=24'b101000010111110100111110;
#1 $display("%b", po);
# 1  pi=24'b111100001011001010111111;
#1 $display("%b", po);
# 1  pi=24'b011111100001100111101000;
#1 $display("%b", po);
# 1  pi=24'b000110011010111111011001;
#1 $display("%b", po);
# 1  pi=24'b111000001100011100101100;
#1 $display("%b", po);
# 1  pi=24'b111000000111011001010010;
#1 $display("%b", po);
# 1  pi=24'b100000011000001000001100;
#1 $display("%b", po);
# 1  pi=24'b100111111101000010000000;
#1 $display("%b", po);
# 1  pi=24'b001011011111110010010101;
#1 $display("%b", po);
# 1  pi=24'b111011011110110110011111;
#1 $display("%b", po);
# 1  pi=24'b110001000000010011110111;
#1 $display("%b", po);
# 1  pi=24'b010001101000000011001010;
#1 $display("%b", po);
# 1  pi=24'b001101101000110100011000;
#1 $display("%b", po);
# 1  pi=24'b001011100010011111010110;
#1 $display("%b", po);
# 1  pi=24'b111010010100001001010100;
#1 $display("%b", po);
# 1  pi=24'b011011110000100010010000;
#1 $display("%b", po);
# 1  pi=24'b110100001101100001000000;
#1 $display("%b", po);
# 1  pi=24'b101001001111110011110010;
#1 $display("%b", po);
# 1  pi=24'b001000010000010110011011;
#1 $display("%b", po);
# 1  pi=24'b101001011010101010100011;
#1 $display("%b", po);
# 1  pi=24'b011111100010111011010011;
#1 $display("%b", po);
# 1  pi=24'b010000101111000100000111;
#1 $display("%b", po);
# 1  pi=24'b111001111000010110010001;
#1 $display("%b", po);
# 1  pi=24'b010110100100010100011101;
#1 $display("%b", po);
# 1  pi=24'b010111101100101110101110;
#1 $display("%b", po);
# 1  pi=24'b111001010111101011111001;
#1 $display("%b", po);
# 1  pi=24'b111010010110110001101000;
#1 $display("%b", po);
# 1  pi=24'b111110000010100110001001;
#1 $display("%b", po);
# 1  pi=24'b111001011111111010010100;
#1 $display("%b", po);
# 1  pi=24'b010110001001111010101100;
#1 $display("%b", po);
# 1  pi=24'b000010011010000101001000;
#1 $display("%b", po);
# 1  pi=24'b100111110010100001000011;
#1 $display("%b", po);
# 1  pi=24'b100000100100000101010111;
#1 $display("%b", po);
# 1  pi=24'b100011001111110101101000;
#1 $display("%b", po);
# 1  pi=24'b000011010110011101101011;
#1 $display("%b", po);
# 1  pi=24'b110000001000101111001111;
#1 $display("%b", po);
# 1  pi=24'b100101001110011101000100;
#1 $display("%b", po);
# 1  pi=24'b110000001001010011101011;
#1 $display("%b", po);
# 1  pi=24'b101100101101000101111101;
#1 $display("%b", po);
# 1  pi=24'b010000111111011100001011;
#1 $display("%b", po);
# 1  pi=24'b110101001000010111000001;
#1 $display("%b", po);
# 1  pi=24'b100000110010111000110011;
#1 $display("%b", po);
end
endmodule

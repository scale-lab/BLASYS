module adder_28(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, po0, po1, po2, po3, po4);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
  output po0, po1, po2, po3, po4;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  assign n9 = pi0 & ~pi4;
  assign n10 = ~pi0 & pi4;
  assign n11 = ~n9 & ~n10;
  assign n12 = pi0 & pi4;
  assign n13 = ~pi1 & ~pi5;
  assign n14 = pi1 & pi5;
  assign n15 = ~n13 & ~n14;
  assign n16 = n12 & ~n15;
  assign n17 = ~n12 & n15;
  assign n18 = ~n16 & ~n17;
  assign n19 = n12 & ~n13;
  assign n20 = ~n14 & ~n19;
  assign n21 = ~pi2 & ~pi6;
  assign n22 = pi2 & pi6;
  assign n23 = ~n21 & ~n22;
  assign n24 = n20 & ~n23;
  assign n25 = ~n20 & n23;
  assign n26 = ~n24 & ~n25;
  assign n27 = ~n20 & ~n21;
  assign n28 = ~n22 & ~n27;
  assign n29 = ~pi3 & ~pi7;
  assign n30 = pi3 & pi7;
  assign n31 = ~n29 & ~n30;
  assign n32 = n28 & ~n31;
  assign n33 = ~n28 & n31;
  assign n34 = ~n32 & ~n33;
  assign n35 = ~n28 & ~n29;
  assign n36 = ~n30 & ~n35;
  assign po0 = n11;
  assign po1 = n18;
  assign po2 = n26;
  assign po3 = n34;
  assign po4 = n36;
endmodule

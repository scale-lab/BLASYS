module adder(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128);
  input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, tpo000, tpo001, tpo002, tpo003, tpo004, tpo005, tpo006, tpo007, tpo008, tpo009, tpo010, tpo011, tpo012, tpo013, tpo014, tpo015, tpo016, tpo017, tpo018, tpo019, tpo020, tpo021, tpo022, tpo023, tpo024, tpo025, tpo026, tpo027, tpo028, tpo029, tpo030, tpo031, tpo032, tpo033, tpo034, tpo035, tpo036, tpo037, tpo038, tpo039, tpo040, tpo041, tpo042, tpo043, tpo044, tpo045, tpo046, tpo047, tpo048, tpo049, tpo050, tpo051, tpo052, tpo053, tpo054, tpo055, tpo056, tpo057, tpo058, tpo059, tpo060, tpo061, tpo062, tpo063, tpo064, tpo065, tpo066, tpo067, tpo068, tpo069, tpo070, tpo071, tpo072, tpo073, tpo074, tpo075, tpo076, tpo077, tpo078, tpo079, tpo080, tpo081, tpo082, tpo083, tpo084, tpo085, tpo086, tpo087, tpo088, tpo089, tpo090, tpo091, tpo092, tpo093, tpo094, tpo095, tpo096, tpo097, tpo098, tpo099, tpo100, tpo101, tpo102, tpo103, tpo104, tpo105, tpo106, tpo107, tpo108, tpo109, tpo110, tpo111, tpo112, tpo113, tpo114, tpo115, tpo116, tpo117, tpo118, tpo119, tpo120, tpo121, tpo122, tpo123, tpo124, tpo125, tpo126, tpo127, tpo128;
  assign po000 = ~tpo000;
  assign po001 = ~tpo001;
  assign po002 = tpo002;
  assign po003 = tpo003;
  assign po004 = tpo004;
  assign po005 = tpo005;
  assign po006 = tpo006;
  assign po007 = tpo007;
  assign po008 = tpo008;
  assign po009 = tpo009;
  assign po010 = tpo010;
  assign po011 = tpo011;
  assign po012 = tpo012;
  assign po013 = tpo013;
  assign po014 = tpo014;
  assign po015 = tpo015;
  assign po016 = tpo016;
  assign po017 = tpo017;
  assign po018 = tpo018;
  assign po019 = tpo019;
  assign po020 = tpo020;
  assign po021 = tpo021;
  assign po022 = tpo022;
  assign po023 = tpo023;
  assign po024 = tpo024;
  assign po025 = tpo025;
  assign po026 = tpo026;
  assign po027 = tpo027;
  assign po028 = tpo028;
  assign po029 = tpo029;
  assign po030 = tpo030;
  assign po031 = tpo031;
  assign po032 = tpo032;
  assign po033 = tpo033;
  assign po034 = tpo034;
  assign po035 = tpo035;
  assign po036 = tpo036;
  assign po037 = tpo037;
  assign po038 = tpo038;
  assign po039 = tpo039;
  assign po040 = tpo040;
  assign po041 = tpo041;
  assign po042 = tpo042;
  assign po043 = tpo043;
  assign po044 = tpo044;
  assign po045 = tpo045;
  assign po046 = tpo046;
  assign po047 = tpo047;
  assign po048 = tpo048;
  assign po049 = tpo049;
  assign po050 = tpo050;
  assign po051 = tpo051;
  assign po052 = tpo052;
  assign po053 = tpo053;
  assign po054 = tpo054;
  assign po055 = tpo055;
  assign po056 = tpo056;
  assign po057 = tpo057;
  assign po058 = tpo058;
  assign po059 = tpo059;
  assign po060 = tpo060;
  assign po061 = tpo061;
  assign po062 = tpo062;
  assign po063 = tpo063;
  assign po064 = tpo064;
  assign po065 = tpo065;
  assign po066 = tpo066;
  assign po067 = tpo067;
  assign po068 = tpo068;
  assign po069 = tpo069;
  assign po070 = tpo070;
  assign po071 = tpo071;
  assign po072 = tpo072;
  assign po073 = tpo073;
  assign po074 = tpo074;
  assign po075 = tpo075;
  assign po076 = tpo076;
  assign po077 = tpo077;
  assign po078 = tpo078;
  assign po079 = tpo079;
  assign po080 = tpo080;
  assign po081 = tpo081;
  assign po082 = tpo082;
  assign po083 = tpo083;
  assign po084 = tpo084;
  assign po085 = tpo085;
  assign po086 = tpo086;
  assign po087 = tpo087;
  assign po088 = tpo088;
  assign po089 = tpo089;
  assign po090 = tpo090;
  assign po091 = tpo091;
  assign po092 = tpo092;
  assign po093 = tpo093;
  assign po094 = tpo094;
  assign po095 = tpo095;
  assign po096 = tpo096;
  assign po097 = tpo097;
  assign po098 = tpo098;
  assign po099 = tpo099;
  assign po100 = tpo100;
  assign po101 = tpo101;
  assign po102 = tpo102;
  assign po103 = tpo103;
  assign po104 = tpo104;
  assign po105 = tpo105;
  assign po106 = tpo106;
  assign po107 = tpo107;
  assign po108 = tpo108;
  assign po109 = tpo109;
  assign po110 = tpo110;
  assign po111 = tpo111;
  assign po112 = tpo112;
  assign po113 = tpo113;
  assign po114 = tpo114;
  assign po115 = tpo115;
  assign po116 = tpo116;
  assign po117 = tpo117;
  assign po118 = tpo118;
  assign po119 = tpo119;
  assign po120 = tpo120;
  assign po121 = tpo121;
  assign po122 = tpo122;
  assign po123 = tpo123;
  assign po124 = tpo124;
  assign po125 = tpo125;
  assign po126 = tpo126;
  assign po127 = tpo127;
  assign po128 = ~tpo128;
  adder_0 U0 ( .pi0( pi115 ), .pi1( pi116 ), .pi2( pi117 ), .pi3( pi243 ), .pi4( pi244 ), .pi5( pi245 ), .pi6( n35 ), .po0( tpo115 ), .po1( tpo116 ), .po2( tpo117 ), .po3( n36 ) );
  adder_1 U1 ( .pi0( pi112 ), .pi1( pi113 ), .pi2( pi114 ), .pi3( pi240 ), .pi4( pi241 ), .pi5( pi242 ), .pi6( n34 ), .po0( tpo112 ), .po1( tpo113 ), .po2( tpo114 ), .po3( n35 ) );
  adder_2 U2 ( .pi0( pi125 ), .pi1( pi126 ), .pi2( pi127 ), .pi3( pi253 ), .pi4( pi254 ), .pi5( pi255 ), .pi6( n38 ), .po0( tpo125 ), .po1( tpo126 ), .po2( tpo127 ), .po3( tpo128 ) );
  adder_3 U3 ( .pi0( pi122 ), .pi1( pi123 ), .pi2( pi124 ), .pi3( pi250 ), .pi4( pi251 ), .pi5( pi252 ), .pi6( n37 ), .po0( tpo122 ), .po1( tpo123 ), .po2( tpo124 ), .po3( n38 ) );
  adder_4 U4 ( .pi0( pi118 ), .pi1( pi119 ), .pi2( pi120 ), .pi3( pi121 ), .pi4( pi246 ), .pi5( pi247 ), .pi6( pi248 ), .pi7( pi249 ), .pi8( n36 ), .po0( tpo118 ), .po1( tpo119 ), .po2( tpo120 ), .po3( tpo121 ), .po4( n37 ) );
  adder_5 U5 ( .pi0( pi106 ), .pi1( pi107 ), .pi2( pi108 ), .pi3( pi234 ), .pi4( pi235 ), .pi5( pi236 ), .pi6( n32 ), .po0( tpo106 ), .po1( tpo107 ), .po2( tpo108 ), .po3( n33 ) );
  adder_6 U6 ( .pi0( pi109 ), .pi1( pi110 ), .pi2( pi111 ), .pi3( pi237 ), .pi4( pi238 ), .pi5( pi239 ), .pi6( n33 ), .po0( tpo109 ), .po1( tpo110 ), .po2( tpo111 ), .po3( n34 ) );
  adder_7 U7 ( .pi0( pi103 ), .pi1( pi104 ), .pi2( pi105 ), .pi3( pi231 ), .pi4( pi232 ), .pi5( pi233 ), .pi6( n31 ), .po0( tpo103 ), .po1( tpo104 ), .po2( tpo105 ), .po3( n32 ) );
  adder_8 U8 ( .pi0( pi096 ), .pi1( pi097 ), .pi2( pi098 ), .pi3( pi224 ), .pi4( pi225 ), .pi5( pi226 ), .pi6( n29 ), .po0( tpo096 ), .po1( tpo097 ), .po2( tpo098 ), .po3( n30 ) );
  adder_9 U9 ( .pi0( pi099 ), .pi1( pi100 ), .pi2( pi101 ), .pi3( pi102 ), .pi4( pi227 ), .pi5( pi228 ), .pi6( pi229 ), .pi7( pi230 ), .pi8( n30 ), .po0( tpo099 ), .po1( tpo100 ), .po2( tpo101 ), .po3( tpo102 ), .po4( n31 ) );
  adder_10 U10 ( .pi0( pi093 ), .pi1( pi094 ), .pi2( pi095 ), .pi3( pi221 ), .pi4( pi222 ), .pi5( pi223 ), .pi6( n28 ), .po0( tpo093 ), .po1( tpo094 ), .po2( tpo095 ), .po3( n29 ) );
  adder_11 U11 ( .pi0( pi090 ), .pi1( pi091 ), .pi2( pi092 ), .pi3( pi218 ), .pi4( pi219 ), .pi5( pi220 ), .pi6( n27 ), .po0( tpo090 ), .po1( tpo091 ), .po2( tpo092 ), .po3( n28 ) );
  adder_12 U12 ( .pi0( pi080 ), .pi1( pi081 ), .pi2( pi082 ), .pi3( pi208 ), .pi4( pi209 ), .pi5( pi210 ), .pi6( n24 ), .po0( tpo080 ), .po1( tpo081 ), .po2( tpo082 ), .po3( n25 ) );
  adder_13 U13 ( .pi0( pi087 ), .pi1( pi088 ), .pi2( pi089 ), .pi3( pi215 ), .pi4( pi216 ), .pi5( pi217 ), .pi6( n26 ), .po0( tpo087 ), .po1( tpo088 ), .po2( tpo089 ), .po3( n27 ) );
  adder_14 U14 ( .pi0( pi083 ), .pi1( pi084 ), .pi2( pi085 ), .pi3( pi086 ), .pi4( pi211 ), .pi5( pi212 ), .pi6( pi213 ), .pi7( pi214 ), .pi8( n25 ), .po0( tpo083 ), .po1( tpo084 ), .po2( tpo085 ), .po3( tpo086 ), .po4( n26 ) );
  adder_15 U15 ( .pi0( pi074 ), .pi1( pi075 ), .pi2( pi076 ), .pi3( pi202 ), .pi4( pi203 ), .pi5( pi204 ), .pi6( n22 ), .po0( tpo074 ), .po1( tpo075 ), .po2( tpo076 ), .po3( n23 ) );
  adder_16 U16 ( .pi0( pi077 ), .pi1( pi078 ), .pi2( pi079 ), .pi3( pi205 ), .pi4( pi206 ), .pi5( pi207 ), .pi6( n23 ), .po0( tpo077 ), .po1( tpo078 ), .po2( tpo079 ), .po3( n24 ) );
  adder_17 U17 ( .pi0( pi071 ), .pi1( pi072 ), .pi2( pi073 ), .pi3( pi199 ), .pi4( pi200 ), .pi5( pi201 ), .pi6( n21 ), .po0( tpo071 ), .po1( tpo072 ), .po2( tpo073 ), .po3( n22 ) );
  adder_18 U18 ( .pi0( pi068 ), .pi1( pi069 ), .pi2( pi070 ), .pi3( pi196 ), .pi4( pi197 ), .pi5( pi198 ), .pi6( n20 ), .po0( tpo068 ), .po1( tpo069 ), .po2( tpo070 ), .po3( n21 ) );
  adder_19 U19 ( .pi0( pi064 ), .pi1( pi065 ), .pi2( pi066 ), .pi3( pi067 ), .pi4( pi192 ), .pi5( pi193 ), .pi6( pi194 ), .pi7( pi195 ), .pi8( n19 ), .po0( tpo064 ), .po1( tpo065 ), .po2( tpo066 ), .po3( tpo067 ), .po4( n20 ) );
  adder_20 U20 ( .pi0( pi016 ), .pi1( pi017 ), .pi2( pi018 ), .pi3( pi144 ), .pi4( pi145 ), .pi5( pi146 ), .pi6( n4 ), .po0( tpo016 ), .po1( tpo017 ), .po2( tpo018 ), .po3( n5 ) );
  adder_21 U21 ( .pi0( pi019 ), .pi1( pi020 ), .pi2( pi021 ), .pi3( pi147 ), .pi4( pi148 ), .pi5( pi149 ), .pi6( n5 ), .po0( tpo019 ), .po1( tpo020 ), .po2( tpo021 ), .po3( n6 ) );
  adder_22 U22 ( .pi0( pi029 ), .pi1( pi030 ), .pi2( pi031 ), .pi3( pi157 ), .pi4( pi158 ), .pi5( pi159 ), .pi6( n8 ), .po0( tpo029 ), .po1( tpo030 ), .po2( tpo031 ), .po3( n9 ) );
  adder_23 U23 ( .pi0( pi022 ), .pi1( pi023 ), .pi2( pi024 ), .pi3( pi025 ), .pi4( pi150 ), .pi5( pi151 ), .pi6( pi152 ), .pi7( pi153 ), .pi8( n6 ), .po0( tpo022 ), .po1( tpo023 ), .po2( tpo024 ), .po3( tpo025 ), .po4( n7 ) );
  adder_24 U24 ( .pi0( pi026 ), .pi1( pi027 ), .pi2( pi028 ), .pi3( pi154 ), .pi4( pi155 ), .pi5( pi156 ), .pi6( n7 ), .po0( tpo026 ), .po1( tpo027 ), .po2( tpo028 ), .po3( n8 ) );
  adder_25 U25 ( .pi0( pi010 ), .pi1( pi011 ), .pi2( pi012 ), .pi3( pi138 ), .pi4( pi139 ), .pi5( pi140 ), .pi6( n2 ), .po0( tpo010 ), .po1( tpo011 ), .po2( tpo012 ), .po3( n3 ) );
  adder_26 U26 ( .pi0( pi013 ), .pi1( pi014 ), .pi2( pi015 ), .pi3( pi141 ), .pi4( pi142 ), .pi5( pi143 ), .pi6( n3 ), .po0( tpo013 ), .po1( tpo014 ), .po2( tpo015 ), .po3( n4 ) );
  adder_27 U27 ( .pi0( pi007 ), .pi1( pi008 ), .pi2( pi009 ), .pi3( pi135 ), .pi4( pi136 ), .pi5( pi137 ), .pi6( n1 ), .po0( tpo007 ), .po1( tpo008 ), .po2( tpo009 ), .po3( n2 ) );
  adder_28 U28 ( .pi0( pi000 ), .pi1( pi001 ), .pi2( pi002 ), .pi3( pi003 ), .pi4( pi128 ), .pi5( pi129 ), .pi6( pi130 ), .pi7( pi131 ), .po0( tpo000 ), .po1( tpo001 ), .po2( tpo002 ), .po3( tpo003 ), .po4( n0 ) );
  adder_29 U29 ( .pi0( pi004 ), .pi1( pi005 ), .pi2( pi006 ), .pi3( pi132 ), .pi4( pi133 ), .pi5( pi134 ), .pi6( n0 ), .po0( tpo004 ), .po1( tpo005 ), .po2( tpo006 ), .po3( n1 ) );
  adder_30 U30 ( .pi0( pi058 ), .pi1( pi059 ), .pi2( pi060 ), .pi3( pi186 ), .pi4( pi187 ), .pi5( pi188 ), .pi6( n17 ), .po0( tpo058 ), .po1( tpo059 ), .po2( tpo060 ), .po3( n18 ) );
  adder_31 U31 ( .pi0( pi061 ), .pi1( pi062 ), .pi2( pi063 ), .pi3( pi189 ), .pi4( pi190 ), .pi5( pi191 ), .pi6( n18 ), .po0( tpo061 ), .po1( tpo062 ), .po2( tpo063 ), .po3( n19 ) );
  adder_32 U32 ( .pi0( pi055 ), .pi1( pi056 ), .pi2( pi057 ), .pi3( pi183 ), .pi4( pi184 ), .pi5( pi185 ), .pi6( n16 ), .po0( tpo055 ), .po1( tpo056 ), .po2( tpo057 ), .po3( n17 ) );
  adder_33 U33 ( .pi0( pi048 ), .pi1( pi049 ), .pi2( pi050 ), .pi3( pi051 ), .pi4( pi176 ), .pi5( pi177 ), .pi6( pi178 ), .pi7( pi179 ), .pi8( n14 ), .po0( tpo048 ), .po1( tpo049 ), .po2( tpo050 ), .po3( tpo051 ), .po4( n15 ) );
  adder_34 U34 ( .pi0( pi052 ), .pi1( pi053 ), .pi2( pi054 ), .pi3( pi180 ), .pi4( pi181 ), .pi5( pi182 ), .pi6( n15 ), .po0( tpo052 ), .po1( tpo053 ), .po2( tpo054 ), .po3( n16 ) );
  adder_35 U35 ( .pi0( pi045 ), .pi1( pi046 ), .pi2( pi047 ), .pi3( pi173 ), .pi4( pi174 ), .pi5( pi175 ), .pi6( n13 ), .po0( tpo045 ), .po1( tpo046 ), .po2( tpo047 ), .po3( n14 ) );
  adder_36 U36 ( .pi0( pi042 ), .pi1( pi043 ), .pi2( pi044 ), .pi3( pi170 ), .pi4( pi171 ), .pi5( pi172 ), .pi6( n12 ), .po0( tpo042 ), .po1( tpo043 ), .po2( tpo044 ), .po3( n13 ) );
  adder_37 U37 ( .pi0( pi032 ), .pi1( pi033 ), .pi2( pi034 ), .pi3( pi160 ), .pi4( pi161 ), .pi5( pi162 ), .pi6( n9 ), .po0( tpo032 ), .po1( tpo033 ), .po2( tpo034 ), .po3( n10 ) );
  adder_38 U38 ( .pi0( pi035 ), .pi1( pi036 ), .pi2( pi037 ), .pi3( pi163 ), .pi4( pi164 ), .pi5( pi165 ), .pi6( n10 ), .po0( tpo035 ), .po1( tpo036 ), .po2( tpo037 ), .po3( n11 ) );
  adder_39 U39 ( .pi0( pi038 ), .pi1( pi039 ), .pi2( pi040 ), .pi3( pi041 ), .pi4( pi166 ), .pi5( pi167 ), .pi6( pi168 ), .pi7( pi169 ), .pi8( n11 ), .po0( tpo038 ), .po1( tpo039 ), .po2( tpo040 ), .po3( tpo041 ), .po4( n12 ) );
endmodule
